(*blackbox*)

module conv_serializer (CLK,SERIAL_OUT,PAR_IN1,PAR_IN2);
    input wire CLK;
    //input RESET;
    output reg SERIAL_OUT;
    input wire PAR_IN1,PAR_IN2;

endmodule