// This is the unpowered netlist.
module lp_tree_serializer (CLK,
    RESET,
    SERIAL_OUT,
    PAR_IN);
 input CLK;
 input RESET;
 output SERIAL_OUT;
 input [15:0] PAR_IN;

 wire \S0.CLK ;
 wire \S0.RESET ;
 wire \S0.SERIAL_OUT ;
 wire \S0.clk_gen[1].clk_gen[0].clks.clk0_o ;
 wire \S0.clk_gen[1].clk_gen[0].clks.clk90_o ;
 wire \S0.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ;
 wire \S0.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ;
 wire \S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ;
 wire \S0.clk_gen[2].clk_gen[0].clks.clk0_o ;
 wire \S0.clk_gen[2].clk_gen[0].clks.clk90_o ;
 wire \S0.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ;
 wire \S0.clk_gen[2].clk_gen[1].clks.clk0_o ;
 wire \S0.clk_gen[2].clk_gen[1].clks.clk90_o ;
 wire \S0.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ;
 wire \S0.stage_gen[1].mux_gen[0].S.PAR_IN1 ;
 wire \S0.stage_gen[1].mux_gen[0].S.PAR_IN2 ;
 wire \S0.stage_gen[1].mux_gen[1].S.PAR_IN1 ;
 wire \S0.stage_gen[1].mux_gen[1].S.PAR_IN2 ;
 wire \S0.stage_gen[1].mux_gen[2].S.PAR_IN1 ;
 wire \S0.stage_gen[1].mux_gen[3].S.PAR_IN1 ;
 wire \S1.CLK ;
 wire \S1.SERIAL_OUT ;
 wire \S1.clk_gen[1].clk_gen[0].clks.clk0_o ;
 wire \S1.clk_gen[1].clk_gen[0].clks.clk90_o ;
 wire \S1.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ;
 wire \S1.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ;
 wire \S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ;
 wire \S1.clk_gen[2].clk_gen[0].clks.clk0_o ;
 wire \S1.clk_gen[2].clk_gen[0].clks.clk90_o ;
 wire \S1.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ;
 wire \S1.clk_gen[2].clk_gen[1].clks.clk0_o ;
 wire \S1.clk_gen[2].clk_gen[1].clks.clk90_o ;
 wire \S1.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ;
 wire \S1.stage_gen[1].mux_gen[0].S.PAR_IN1 ;
 wire \S1.stage_gen[1].mux_gen[0].S.PAR_IN2 ;
 wire \S1.stage_gen[1].mux_gen[1].S.PAR_IN1 ;
 wire \S1.stage_gen[1].mux_gen[2].S.PAR_IN1 ;
 wire \S1.stage_gen[1].mux_gen[3].S.PAR_IN1 ;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire \clkdiv0.hold_rsts[0] ;
 wire \clkdiv0.hold_rsts[1] ;
 wire clknet_0_CLK;
 wire clknet_1_0__leaf_CLK;
 wire clknet_1_1__leaf_CLK;
 wire \last_stage.PAR_IN1 ;
 wire \last_stage.PAR_IN2 ;
 wire \last_stage_inputs[0] ;
 wire \last_stage_inputs[1] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__nand2_1 _078_ (.A(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _079_ (.A(\S1.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S1.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _080_ (.A(\S1.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ),
    .B(\S1.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _081_ (.A(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_015_));
 sky130_fd_sc_hd__nand2_1 _082_ (.A(\S0.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S0.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _083_ (.A(\S0.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ),
    .B(\S0.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _084_ (.A(\clkdiv0.hold_rsts[0] ),
    .B(\S1.CLK ),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _085_ (.A(net12),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _086_ (.A(\S0.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _087_ (.A(_065_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _088_ (.A(\S0.stage_gen[1].mux_gen[2].S.PAR_IN1 ),
    .Y(_068_));
 sky130_fd_sc_hd__nand2_1 _089_ (.A(_068_),
    .B(\S0.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .Y(_069_));
 sky130_fd_sc_hd__nand3_1 _090_ (.A(_067_),
    .B(_069_),
    .C(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _091_ (.A(net14),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _092_ (.A(\S0.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_072_));
 sky130_fd_sc_hd__nand2_1 _093_ (.A(_071_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _094_ (.A(\S0.stage_gen[1].mux_gen[3].S.PAR_IN1 ),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _095_ (.A(_074_),
    .B(\S0.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_075_));
 sky130_fd_sc_hd__clkinv_4 _096_ (.A(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_001_));
 sky130_fd_sc_hd__nand3_1 _097_ (.A(_073_),
    .B(_075_),
    .C(_001_),
    .Y(_076_));
 sky130_fd_sc_hd__nand2_1 _098_ (.A(_070_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _099_ (.A(\S0.CLK ),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _100_ (.A(_077_),
    .B(_003_),
    .Y(_027_));
 sky130_fd_sc_hd__nand2b_1 _101_ (.A_N(\S0.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .B(\S0.stage_gen[1].mux_gen[1].S.PAR_IN2 ),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _102_ (.A(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_1 _103_ (.A(\S0.stage_gen[1].mux_gen[1].S.PAR_IN1 ),
    .B(\S0.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .Y(_029_));
 sky130_fd_sc_hd__nand3_1 _104_ (.A(_028_),
    .B(_002_),
    .C(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _105_ (.A(\S0.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _106_ (.A(_031_),
    .B(\S0.stage_gen[1].mux_gen[0].S.PAR_IN2 ),
    .Y(_032_));
 sky130_fd_sc_hd__nand2_1 _107_ (.A(\S0.stage_gen[1].mux_gen[0].S.PAR_IN1 ),
    .B(\S0.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .Y(_033_));
 sky130_fd_sc_hd__nand3_1 _108_ (.A(_032_),
    .B(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .C(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__nand3_1 _109_ (.A(_030_),
    .B(_034_),
    .C(\S0.CLK ),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _110_ (.A(_027_),
    .B(_035_),
    .Y(\S0.SERIAL_OUT ));
 sky130_fd_sc_hd__inv_2 _111_ (.A(net5),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _112_ (.A(\S1.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _113_ (.A(_036_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _114_ (.A(\S1.stage_gen[1].mux_gen[2].S.PAR_IN1 ),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _115_ (.A(_039_),
    .B(\S1.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .Y(_040_));
 sky130_fd_sc_hd__nand3_1 _116_ (.A(_038_),
    .B(_040_),
    .C(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(net7),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _118_ (.A(\S1.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _119_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _120_ (.A(\S1.stage_gen[1].mux_gen[3].S.PAR_IN1 ),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_1 _121_ (.A(_045_),
    .B(\S1.clk_gen[2].clk_gen[1].clks.clk90_o ),
    .Y(_046_));
 sky130_fd_sc_hd__clkinv_4 _122_ (.A(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .Y(_004_));
 sky130_fd_sc_hd__nand3_1 _123_ (.A(_044_),
    .B(_046_),
    .C(_004_),
    .Y(_047_));
 sky130_fd_sc_hd__nand2_1 _124_ (.A(_041_),
    .B(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _125_ (.A(\S1.CLK ),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _126_ (.A(_048_),
    .B(_006_),
    .Y(_049_));
 sky130_fd_sc_hd__nand2b_1 _127_ (.A_N(\S1.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .B(net3),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _128_ (.A(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _129_ (.A(\S1.stage_gen[1].mux_gen[1].S.PAR_IN1 ),
    .B(\S1.clk_gen[2].clk_gen[0].clks.clk90_o ),
    .Y(_051_));
 sky130_fd_sc_hd__nand3_1 _130_ (.A(_050_),
    .B(_005_),
    .C(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _131_ (.A(\S1.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .Y(_053_));
 sky130_fd_sc_hd__nand2_1 _132_ (.A(_053_),
    .B(\S1.stage_gen[1].mux_gen[0].S.PAR_IN2 ),
    .Y(_054_));
 sky130_fd_sc_hd__nand2_1 _133_ (.A(\S1.stage_gen[1].mux_gen[0].S.PAR_IN1 ),
    .B(\S1.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .Y(_055_));
 sky130_fd_sc_hd__nand3_1 _134_ (.A(_054_),
    .B(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .C(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__nand3_1 _135_ (.A(_052_),
    .B(_056_),
    .C(\S1.CLK ),
    .Y(_057_));
 sky130_fd_sc_hd__nand2_1 _136_ (.A(_049_),
    .B(_057_),
    .Y(\S1.SERIAL_OUT ));
 sky130_fd_sc_hd__mux2_4 _137_ (.A0(\last_stage.PAR_IN2 ),
    .A1(\last_stage.PAR_IN1 ),
    .S(clknet_1_0__leaf_CLK),
    .X(_058_));
 sky130_fd_sc_hd__buf_6 _138_ (.A(_058_),
    .X(net18));
 sky130_fd_sc_hd__nand2_1 _139_ (.A(\S0.CLK ),
    .B(net17),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _140__1 (.A(clknet_1_1__leaf_CLK),
    .Y(net19));
 sky130_fd_sc_hd__nand2_1 _141_ (.A(\S0.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .B(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Y(_010_));
 sky130_fd_sc_hd__nand2_1 _142_ (.A(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S0.RESET ),
    .Y(_059_));
 sky130_fd_sc_hd__clkinv_2 _143_ (.A(_059_),
    .Y(_011_));
 sky130_fd_sc_hd__nand2_1 _144_ (.A(\S0.RESET ),
    .B(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ),
    .Y(_060_));
 sky130_fd_sc_hd__clkinv_2 _145_ (.A(_060_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _146_ (.A(\S0.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .B(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _147_ (.A(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .B(\S0.RESET ),
    .Y(_016_));
 sky130_fd_sc_hd__nand2_1 _148_ (.A(\clkdiv0.hold_rsts[0] ),
    .B(net17),
    .Y(_061_));
 sky130_fd_sc_hd__clkinv_2 _149_ (.A(_061_),
    .Y(_017_));
 sky130_fd_sc_hd__nand2_1 _150_ (.A(net17),
    .B(\clkdiv0.hold_rsts[1] ),
    .Y(_062_));
 sky130_fd_sc_hd__clkinv_2 _151_ (.A(_062_),
    .Y(_018_));
 sky130_fd_sc_hd__nand2_1 _152_ (.A(\S1.clk_gen[2].clk_gen[1].clks.clk0_o ),
    .B(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Y(_020_));
 sky130_fd_sc_hd__nand2_1 _153_ (.A(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ),
    .B(\S0.RESET ),
    .Y(_063_));
 sky130_fd_sc_hd__clkinv_2 _154_ (.A(_063_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _155_ (.A(\S0.RESET ),
    .B(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ),
    .Y(_064_));
 sky130_fd_sc_hd__clkinv_2 _156_ (.A(_064_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _157_ (.A(\S1.clk_gen[2].clk_gen[0].clks.clk0_o ),
    .B(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _158_ (.A(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .B(\S0.RESET ),
    .Y(_026_));
 sky130_fd_sc_hd__dlxtp_1 _159_ (.D(\S0.SERIAL_OUT ),
    .GATE(clknet_1_0__leaf_CLK),
    .Q(\last_stage_inputs[0] ));
 sky130_fd_sc_hd__dlxtn_1 _160_ (.D(\S1.SERIAL_OUT ),
    .GATE_N(clknet_1_0__leaf_CLK),
    .Q(\last_stage_inputs[1] ));
 sky130_fd_sc_hd__dlxtn_1 _161_ (.D(\last_stage_inputs[0] ),
    .GATE_N(clknet_1_0__leaf_CLK),
    .Q(\last_stage.PAR_IN1 ));
 sky130_fd_sc_hd__dlxtp_1 _162_ (.D(\last_stage_inputs[1] ),
    .GATE(clknet_1_0__leaf_CLK),
    .Q(\last_stage.PAR_IN2 ));
 sky130_fd_sc_hd__dlxtn_1 _163_ (.D(net8),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S0.stage_gen[1].mux_gen[0].S.PAR_IN2 ));
 sky130_fd_sc_hd__dlxtn_1 _164_ (.D(net10),
    .GATE_N(clknet_1_0__leaf_CLK),
    .Q(\S0.stage_gen[1].mux_gen[1].S.PAR_IN2 ));
 sky130_fd_sc_hd__dlxtn_1 _165_ (.D(net11),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S0.stage_gen[1].mux_gen[2].S.PAR_IN1 ));
 sky130_fd_sc_hd__dlxtn_1 _166_ (.D(net13),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S0.stage_gen[1].mux_gen[3].S.PAR_IN1 ));
 sky130_fd_sc_hd__dlxtn_1 _167_ (.D(net16),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S1.stage_gen[1].mux_gen[0].S.PAR_IN2 ));
 sky130_fd_sc_hd__dlxtn_1 _168_ (.D(net2),
    .GATE_N(clknet_1_0__leaf_CLK),
    .Q(\S1.stage_gen[1].mux_gen[1].S.PAR_IN1 ));
 sky130_fd_sc_hd__dlxtn_1 _169_ (.D(net4),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S1.stage_gen[1].mux_gen[2].S.PAR_IN1 ));
 sky130_fd_sc_hd__dlxtn_1 _170_ (.D(net6),
    .GATE_N(clknet_1_1__leaf_CLK),
    .Q(\S1.stage_gen[1].mux_gen[3].S.PAR_IN1 ));
 sky130_fd_sc_hd__dfxtp_1 _171_ (.CLK(clknet_1_0__leaf_CLK),
    .D(net1),
    .Q(\S0.stage_gen[1].mux_gen[0].S.PAR_IN1 ));
 sky130_fd_sc_hd__dfxtp_1 _172_ (.CLK(clknet_1_0__leaf_CLK),
    .D(net9),
    .Q(\S0.stage_gen[1].mux_gen[1].S.PAR_IN1 ));
 sky130_fd_sc_hd__dfxtp_1 _173_ (.CLK(clknet_1_0__leaf_CLK),
    .D(net15),
    .Q(\S1.stage_gen[1].mux_gen[0].S.PAR_IN1 ));
 sky130_fd_sc_hd__dfxtp_2 _174_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_007_),
    .Q(\S0.CLK ));
 sky130_fd_sc_hd__dfxtp_1 _175_ (.CLK(net19),
    .D(_008_),
    .Q(\S1.CLK ));
 sky130_fd_sc_hd__dfxtp_1 _176_ (.CLK(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .D(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Q(\S1.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _177_ (.CLK(_001_),
    .D(_009_),
    .Q(\S0.clk_gen[2].clk_gen[1].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _178_ (.CLK(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .D(_010_),
    .Q(\S0.clk_gen[2].clk_gen[1].clks.clk0_o ));
 sky130_fd_sc_hd__dfxtp_1 _179_ (.CLK(\S0.CLK ),
    .D(_011_),
    .Q(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ));
 sky130_fd_sc_hd__dfxtp_1 _180_ (.CLK(\S0.CLK ),
    .D(_012_),
    .Q(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ));
 sky130_fd_sc_hd__dfxtp_1 _181_ (.CLK(_002_),
    .D(_013_),
    .Q(\S0.clk_gen[2].clk_gen[0].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _182_ (.CLK(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .D(_014_),
    .Q(\S0.clk_gen[2].clk_gen[0].clks.clk0_o ));
 sky130_fd_sc_hd__dfxtp_1 _183_ (.CLK(_003_),
    .D(_015_),
    .Q(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _184_ (.CLK(\S0.CLK ),
    .D(_016_),
    .Q(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ));
 sky130_fd_sc_hd__dfxtp_1 _185_ (.CLK(\S0.CLK ),
    .D(\S0.RESET ),
    .Q(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _186_ (.CLK(\S0.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .D(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Q(\S0.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _187_ (.CLK(\S0.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .D(\S0.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Q(\S0.clk_gen[2].clk_gen[1].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _188_ (.CLK(\S1.CLK ),
    .D(\S0.RESET ),
    .Q(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _189_ (.CLK(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .D(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ),
    .Q(\S1.clk_gen[2].clk_gen[0].clks.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _190_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_017_),
    .Q(\clkdiv0.hold_rsts[1] ));
 sky130_fd_sc_hd__dfxtp_2 _191_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_018_),
    .Q(\S0.RESET ));
 sky130_fd_sc_hd__dfxtp_1 _192_ (.CLK(_004_),
    .D(_019_),
    .Q(\S1.clk_gen[2].clk_gen[1].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _193_ (.CLK(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ),
    .D(_020_),
    .Q(\S1.clk_gen[2].clk_gen[1].clks.clk0_o ));
 sky130_fd_sc_hd__dfxtp_1 _194_ (.CLK(\S1.CLK ),
    .D(_021_),
    .Q(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[1] ));
 sky130_fd_sc_hd__dfxtp_1 _195_ (.CLK(\S1.CLK ),
    .D(_022_),
    .Q(\S1.clk_gen[1].clk_gen[0].clks.hold_rsts[2] ));
 sky130_fd_sc_hd__dfxtp_1 _196_ (.CLK(_005_),
    .D(_023_),
    .Q(\S1.clk_gen[2].clk_gen[0].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _197_ (.CLK(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ),
    .D(_024_),
    .Q(\S1.clk_gen[2].clk_gen[0].clks.clk0_o ));
 sky130_fd_sc_hd__dfxtp_1 _198_ (.CLK(clknet_1_1__leaf_CLK),
    .D(net17),
    .Q(\clkdiv0.hold_rsts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _199_ (.CLK(_006_),
    .D(_025_),
    .Q(\S1.clk_gen[1].clk_gen[0].clks.clk90_o ));
 sky130_fd_sc_hd__dfxtp_1 _200_ (.CLK(\S1.CLK ),
    .D(_026_),
    .Q(\S1.clk_gen[1].clk_gen[0].clks.clk0_o ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(PAR_IN[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(PAR_IN[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(PAR_IN[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(PAR_IN[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(PAR_IN[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(PAR_IN[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(PAR_IN[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(PAR_IN[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(RESET),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(PAR_IN[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(PAR_IN[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(PAR_IN[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(PAR_IN[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(PAR_IN[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(PAR_IN[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(PAR_IN[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(PAR_IN[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 output18 (.A(net18),
    .X(SERIAL_OUT));
endmodule

