// This is the unpowered netlist.
module serializer_unit_cell (CLK,
    COMPLETE,
    INTERNAL_FINISH,
    READY,
    RESET,
    SERIAL_OUT,
    COUNT,
    PAR_IN1,
    PAR_IN2,
    PAR_IN3,
    PAR_IN4,
    PAR_IN5,
    PAR_IN6,
    PAR_IN7,
    PAR_IN8,
    SAMPLE_COUNT);
 input CLK;
 output COMPLETE;
 output INTERNAL_FINISH;
 input READY;
 input RESET;
 output SERIAL_OUT;
 output [5:0] COUNT;
 input [31:0] PAR_IN1;
 input [31:0] PAR_IN2;
 input [31:0] PAR_IN3;
 input [31:0] PAR_IN4;
 input [31:0] PAR_IN5;
 input [31:0] PAR_IN6;
 input [31:0] PAR_IN7;
 input [31:0] PAR_IN8;
 output [3:0] SAMPLE_COUNT;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire clknet_0_CLK;
 wire clknet_1_0__leaf_CLK;
 wire clknet_1_1__leaf_CLK;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net270));
 sky130_fd_sc_hd__fill_2 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__nand2_2 _0676_ (.A(net261),
    .B(net260),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0013_),
    .Y(_0014_));
 sky130_fd_sc_hd__and3_1 _0678_ (.A(_0014_),
    .B(net263),
    .C(net262),
    .X(_0015_));
 sky130_fd_sc_hd__a21o_1 _0679_ (.A1(_0015_),
    .A2(net264),
    .B1(net265),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_2 _0680_ (.A(net267),
    .B(net268),
    .Y(_0017_));
 sky130_fd_sc_hd__clkinv_2 _0681_ (.A(net272),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _0682_ (.A(_0018_),
    .B(net269),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_1 _0683_ (.A(_0017_),
    .B(_0019_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_2 _0684_ (.A(_0020_),
    .X(_0021_));
 sky130_fd_sc_hd__a21bo_1 _0685_ (.A1(net272),
    .A2(net266),
    .B1_N(net257),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _0686_ (.A(net259),
    .B(_0022_),
    .Y(_0023_));
 sky130_fd_sc_hd__and3_1 _0687_ (.A(_0016_),
    .B(_0021_),
    .C(_0023_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0024_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(_0023_),
    .Y(_0025_));
 sky130_fd_sc_hd__or3_1 _0690_ (.A(net272),
    .B(_0025_),
    .C(_0016_),
    .X(_0026_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(net259),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_1 _0692_ (.A(_0027_),
    .B(_0022_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand2_2 _0694_ (.A(_0026_),
    .B(_0029_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(net267),
    .Y(_0031_));
 sky130_fd_sc_hd__nor2_1 _0696_ (.A(_0018_),
    .B(_0025_),
    .Y(_0032_));
 sky130_fd_sc_hd__a31o_1 _0697_ (.A1(_0016_),
    .A2(_0031_),
    .A3(_0023_),
    .B1(_0032_),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _0698_ (.A1(_0030_),
    .A2(net267),
    .B1(_0033_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_2 _0699_ (.A(net268),
    .B(_0031_),
    .Y(_0034_));
 sky130_fd_sc_hd__buf_6 _0700_ (.A(_0034_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_6 _0701_ (.A(_0035_),
    .X(_0036_));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(net268),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _0703_ (.A(net267),
    .B(_0037_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_6 _0704_ (.A(_0038_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_6 _0705_ (.A(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__o211a_1 _0706_ (.A1(_0036_),
    .A2(_0040_),
    .B1(net257),
    .C1(_0018_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(_0041_),
    .A1(net268),
    .S(_0030_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_1 _0708_ (.A(_0042_),
    .X(_0002_));
 sky130_fd_sc_hd__a21oi_1 _0709_ (.A1(net257),
    .A2(_0018_),
    .B1(_0030_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(net269),
    .Y(_0044_));
 sky130_fd_sc_hd__nor3_1 _0711_ (.A(_0044_),
    .B(_0017_),
    .C(_0030_),
    .Y(_0045_));
 sky130_fd_sc_hd__o21ai_1 _0712_ (.A1(_0017_),
    .A2(_0030_),
    .B1(_0044_),
    .Y(_0046_));
 sky130_fd_sc_hd__nor3b_1 _0713_ (.A(_0043_),
    .B(_0045_),
    .C_N(_0046_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ba_1 _0714_ (.A1(net272),
    .A2(_0045_),
    .B1_N(_0022_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0047_),
    .X(_0004_));
 sky130_fd_sc_hd__nor2_1 _0716_ (.A(net272),
    .B(_0044_),
    .Y(_0048_));
 sky130_fd_sc_hd__buf_4 _0717_ (.A(_0048_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_4 _0718_ (.A(_0049_),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_4 _0719_ (.A(_0038_),
    .X(_0051_));
 sky130_fd_sc_hd__nand3_1 _0720_ (.A(_0050_),
    .B(_0051_),
    .C(net202),
    .Y(_0052_));
 sky130_fd_sc_hd__clkinv_4 _0721_ (.A(_0017_),
    .Y(_0053_));
 sky130_fd_sc_hd__buf_2 _0722_ (.A(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__nor2_1 _0723_ (.A(net269),
    .B(net272),
    .Y(_0055_));
 sky130_fd_sc_hd__clkbuf_2 _0724_ (.A(_0055_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_2 _0725_ (.A(_0056_),
    .X(_0057_));
 sky130_fd_sc_hd__nand3_1 _0726_ (.A(_0054_),
    .B(_0057_),
    .C(net106),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _0727_ (.A(_0052_),
    .B(_0058_),
    .Y(_0059_));
 sky130_fd_sc_hd__clkbuf_4 _0728_ (.A(_0049_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_6 _0729_ (.A(_0035_),
    .X(_0061_));
 sky130_fd_sc_hd__nand3_1 _0730_ (.A(_0060_),
    .B(_0061_),
    .C(net170),
    .Y(_0062_));
 sky130_fd_sc_hd__buf_2 _0731_ (.A(_0055_),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_4 _0732_ (.A(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__nand3_1 _0733_ (.A(_0036_),
    .B(net42),
    .C(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__nand2_1 _0734_ (.A(_0062_),
    .B(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__nor2_1 _0735_ (.A(_0059_),
    .B(_0066_),
    .Y(_0067_));
 sky130_fd_sc_hd__buf_4 _0736_ (.A(_0049_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_2 _0737_ (.A(_0053_),
    .X(_0069_));
 sky130_fd_sc_hd__nand3_1 _0738_ (.A(_0068_),
    .B(_0069_),
    .C(net234),
    .Y(_0070_));
 sky130_fd_sc_hd__clkbuf_4 _0739_ (.A(_0056_),
    .X(_0071_));
 sky130_fd_sc_hd__nand3_1 _0740_ (.A(_0051_),
    .B(net74),
    .C(_0071_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _0741_ (.A(_0070_),
    .B(_0072_),
    .Y(_0073_));
 sky130_fd_sc_hd__o21bai_4 _0742_ (.A1(net267),
    .A2(net268),
    .B1_N(net272),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(_0074_),
    .B(_0019_),
    .Y(_0075_));
 sky130_fd_sc_hd__clkbuf_4 _0744_ (.A(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _0745_ (.A(_0074_),
    .B(net138),
    .Y(_0077_));
 sky130_fd_sc_hd__nand2_1 _0746_ (.A(_0076_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor2_1 _0747_ (.A(_0073_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _0748_ (.A(_0067_),
    .B(_0079_),
    .Y(_0080_));
 sky130_fd_sc_hd__buf_2 _0749_ (.A(_0075_),
    .X(_0081_));
 sky130_fd_sc_hd__or2_1 _0750_ (.A(net10),
    .B(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _0751_ (.A(_0080_),
    .B(_0082_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(net261),
    .Y(_0084_));
 sky130_fd_sc_hd__nor2_1 _0753_ (.A(net260),
    .B(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__a21oi_1 _0754_ (.A1(_0083_),
    .A2(_0085_),
    .B1(net262),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_1 _0755_ (.A(_0021_),
    .B(net232),
    .Y(_0087_));
 sky130_fd_sc_hd__buf_2 _0756_ (.A(_0063_),
    .X(_0088_));
 sky130_fd_sc_hd__nand3_1 _0757_ (.A(_0036_),
    .B(net40),
    .C(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0087_),
    .B(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(net104),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_4 _0760_ (.A(_0053_),
    .B(_0063_),
    .Y(_0092_));
 sky130_fd_sc_hd__buf_4 _0761_ (.A(_0048_),
    .X(_0093_));
 sky130_fd_sc_hd__buf_4 _0762_ (.A(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__nand3_1 _0763_ (.A(_0094_),
    .B(_0036_),
    .C(net168),
    .Y(_0095_));
 sky130_fd_sc_hd__o21ai_1 _0764_ (.A1(_0091_),
    .A2(_0092_),
    .B1(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nor2_1 _0765_ (.A(_0090_),
    .B(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__buf_2 _0766_ (.A(_0049_),
    .X(_0098_));
 sky130_fd_sc_hd__buf_6 _0767_ (.A(_0039_),
    .X(_0099_));
 sky130_fd_sc_hd__nand3_1 _0768_ (.A(_0098_),
    .B(_0099_),
    .C(net200),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _0769_ (.A(_0074_),
    .B(net136),
    .Y(_0101_));
 sky130_fd_sc_hd__nand2_1 _0770_ (.A(_0100_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(net72),
    .Y(_0103_));
 sky130_fd_sc_hd__nand2_1 _0772_ (.A(_0039_),
    .B(_0063_),
    .Y(_0104_));
 sky130_fd_sc_hd__buf_2 _0773_ (.A(_0075_),
    .X(_0105_));
 sky130_fd_sc_hd__o21ai_1 _0774_ (.A1(_0103_),
    .A2(_0104_),
    .B1(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__nor2_1 _0775_ (.A(_0102_),
    .B(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _0776_ (.A(_0097_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__buf_2 _0777_ (.A(_0075_),
    .X(_0109_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(net260),
    .Y(_0110_));
 sky130_fd_sc_hd__buf_2 _0779_ (.A(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__o21a_1 _0780_ (.A1(net8),
    .A2(_0109_),
    .B1(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(_0108_),
    .B(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__buf_4 _0782_ (.A(_0049_),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_4 _0783_ (.A(net267),
    .B(net268),
    .Y(_0115_));
 sky130_fd_sc_hd__clkbuf_4 _0784_ (.A(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__nand3_1 _0785_ (.A(_0114_),
    .B(net137),
    .C(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__buf_2 _0786_ (.A(_0056_),
    .X(_0118_));
 sky130_fd_sc_hd__nand3_1 _0787_ (.A(_0054_),
    .B(_0118_),
    .C(net105),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_1 _0788_ (.A(_0117_),
    .B(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand3_1 _0789_ (.A(_0094_),
    .B(_0040_),
    .C(net201),
    .Y(_0121_));
 sky130_fd_sc_hd__buf_6 _0790_ (.A(_0035_),
    .X(_0122_));
 sky130_fd_sc_hd__nand3_1 _0791_ (.A(_0098_),
    .B(_0122_),
    .C(net169),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _0792_ (.A(_0121_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor2_1 _0793_ (.A(_0120_),
    .B(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__buf_6 _0794_ (.A(_0035_),
    .X(_0126_));
 sky130_fd_sc_hd__buf_2 _0795_ (.A(_0056_),
    .X(_0127_));
 sky130_fd_sc_hd__nand3_1 _0796_ (.A(_0126_),
    .B(net41),
    .C(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__buf_2 _0797_ (.A(_0056_),
    .X(_0129_));
 sky130_fd_sc_hd__nand3_1 _0798_ (.A(_0051_),
    .B(net73),
    .C(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _0799_ (.A(_0128_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__clkbuf_4 _0800_ (.A(_0020_),
    .X(_0132_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0132_),
    .B(net233),
    .Y(_0133_));
 sky130_fd_sc_hd__buf_2 _0802_ (.A(_0075_),
    .X(_0134_));
 sky130_fd_sc_hd__nand2_1 _0803_ (.A(_0133_),
    .B(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__nor2_1 _0804_ (.A(_0131_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(_0125_),
    .B(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__buf_2 _0806_ (.A(net260),
    .X(_0138_));
 sky130_fd_sc_hd__o21a_1 _0807_ (.A1(net9),
    .A2(_0105_),
    .B1(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _0808_ (.A(_0137_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__buf_2 _0809_ (.A(_0084_),
    .X(_0141_));
 sky130_fd_sc_hd__nand3_1 _0810_ (.A(_0113_),
    .B(_0140_),
    .C(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(net107),
    .Y(_0143_));
 sky130_fd_sc_hd__buf_2 _0812_ (.A(_0075_),
    .X(_0144_));
 sky130_fd_sc_hd__o21ai_1 _0813_ (.A1(_0143_),
    .A2(_0092_),
    .B1(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(net43),
    .Y(_0146_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(_0034_),
    .B(_0056_),
    .Y(_0147_));
 sky130_fd_sc_hd__clkbuf_4 _0816_ (.A(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(_0021_),
    .B(net235),
    .Y(_0149_));
 sky130_fd_sc_hd__o21ai_1 _0818_ (.A1(_0146_),
    .A2(_0148_),
    .B1(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _0819_ (.A(_0145_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand3_1 _0820_ (.A(_0098_),
    .B(_0122_),
    .C(net171),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(_0074_),
    .B(net139),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _0822_ (.A(_0152_),
    .B(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(net203),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _0824_ (.A(_0048_),
    .B(_0038_),
    .Y(_0156_));
 sky130_fd_sc_hd__buf_2 _0825_ (.A(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__nand3_1 _0826_ (.A(_0040_),
    .B(net75),
    .C(_0088_),
    .Y(_0158_));
 sky130_fd_sc_hd__o21ai_1 _0827_ (.A1(_0155_),
    .A2(_0157_),
    .B1(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _0828_ (.A(_0154_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _0829_ (.A(_0151_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__o21ai_1 _0830_ (.A1(net11),
    .A2(_0109_),
    .B1(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _0831_ (.A(_0162_),
    .B(_0014_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand3_1 _0832_ (.A(_0086_),
    .B(_0142_),
    .C(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(net263),
    .Y(_0165_));
 sky130_fd_sc_hd__nand3_1 _0834_ (.A(_0060_),
    .B(_0061_),
    .C(net176),
    .Y(_0166_));
 sky130_fd_sc_hd__nand3_1 _0835_ (.A(_0040_),
    .B(net80),
    .C(_0064_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(_0166_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(net208),
    .Y(_0169_));
 sky130_fd_sc_hd__clkbuf_4 _0838_ (.A(_0053_),
    .X(_0170_));
 sky130_fd_sc_hd__nand3_1 _0839_ (.A(_0170_),
    .B(_0088_),
    .C(net112),
    .Y(_0171_));
 sky130_fd_sc_hd__o21ai_1 _0840_ (.A1(_0169_),
    .A2(_0157_),
    .B1(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nor2_1 _0841_ (.A(_0168_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__nand3_1 _0842_ (.A(_0122_),
    .B(net48),
    .C(_0118_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _0843_ (.A(_0076_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _0844_ (.A(_0021_),
    .B(net240),
    .Y(_0176_));
 sky130_fd_sc_hd__nand2_1 _0845_ (.A(_0074_),
    .B(net144),
    .Y(_0177_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0175_),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_1 _0848_ (.A(_0173_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__o21a_1 _0849_ (.A1(net16),
    .A2(_0109_),
    .B1(_0138_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _0850_ (.A(_0180_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__buf_6 _0851_ (.A(_0035_),
    .X(_0183_));
 sky130_fd_sc_hd__nand3_1 _0852_ (.A(_0050_),
    .B(_0183_),
    .C(net175),
    .Y(_0184_));
 sky130_fd_sc_hd__nand3_1 _0853_ (.A(_0054_),
    .B(_0127_),
    .C(net111),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _0854_ (.A(_0184_),
    .B(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__buf_6 _0855_ (.A(_0039_),
    .X(_0187_));
 sky130_fd_sc_hd__nand3_1 _0856_ (.A(_0094_),
    .B(_0187_),
    .C(net207),
    .Y(_0188_));
 sky130_fd_sc_hd__nand2_1 _0857_ (.A(_0188_),
    .B(_0076_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _0858_ (.A(_0186_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__buf_2 _0859_ (.A(_0053_),
    .X(_0191_));
 sky130_fd_sc_hd__nand3_1 _0860_ (.A(_0068_),
    .B(_0191_),
    .C(net239),
    .Y(_0192_));
 sky130_fd_sc_hd__nand3_1 _0861_ (.A(_0051_),
    .B(net79),
    .C(_0071_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _0862_ (.A(_0192_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand3_1 _0863_ (.A(_0036_),
    .B(net47),
    .C(_0064_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand3_1 _0864_ (.A(_0050_),
    .B(net143),
    .C(_0116_),
    .Y(_0196_));
 sky130_fd_sc_hd__nand2_1 _0865_ (.A(_0195_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _0866_ (.A(_0194_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(_0190_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__o21a_1 _0868_ (.A1(net15),
    .A2(_0105_),
    .B1(_0111_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _0869_ (.A(_0199_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand3_1 _0870_ (.A(_0182_),
    .B(_0201_),
    .C(net261),
    .Y(_0202_));
 sky130_fd_sc_hd__buf_2 _0871_ (.A(_0038_),
    .X(_0203_));
 sky130_fd_sc_hd__nand3_1 _0872_ (.A(_0203_),
    .B(net78),
    .C(_0057_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _0873_ (.A(_0134_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand3_1 _0874_ (.A(_0094_),
    .B(_0187_),
    .C(net206),
    .Y(_0206_));
 sky130_fd_sc_hd__nand3_1 _0875_ (.A(_0114_),
    .B(net142),
    .C(_0116_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _0876_ (.A(_0206_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(_0205_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand3_1 _0878_ (.A(_0068_),
    .B(_0191_),
    .C(net238),
    .Y(_0210_));
 sky130_fd_sc_hd__nand3_1 _0879_ (.A(_0183_),
    .B(net46),
    .C(_0071_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _0880_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand3_1 _0881_ (.A(_0114_),
    .B(_0126_),
    .C(net174),
    .Y(_0213_));
 sky130_fd_sc_hd__buf_2 _0882_ (.A(_0063_),
    .X(_0214_));
 sky130_fd_sc_hd__nand3_1 _0883_ (.A(_0170_),
    .B(_0214_),
    .C(net110),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0213_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor2_1 _0885_ (.A(_0212_),
    .B(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0209_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__o21a_1 _0887_ (.A1(net14),
    .A2(_0144_),
    .B1(_0138_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_1 _0888_ (.A(_0218_),
    .B(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand3_1 _0889_ (.A(_0183_),
    .B(net45),
    .C(_0129_),
    .Y(_0221_));
 sky130_fd_sc_hd__buf_4 _0890_ (.A(_0049_),
    .X(_0222_));
 sky130_fd_sc_hd__buf_2 _0891_ (.A(_0115_),
    .X(_0223_));
 sky130_fd_sc_hd__nand3_1 _0892_ (.A(_0222_),
    .B(net141),
    .C(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _0893_ (.A(_0221_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand3_1 _0894_ (.A(_0114_),
    .B(_0203_),
    .C(net205),
    .Y(_0226_));
 sky130_fd_sc_hd__nand3_1 _0895_ (.A(_0068_),
    .B(_0183_),
    .C(net173),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _0896_ (.A(_0226_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0225_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand3_1 _0898_ (.A(_0222_),
    .B(_0053_),
    .C(net237),
    .Y(_0230_));
 sky130_fd_sc_hd__buf_2 _0899_ (.A(_0056_),
    .X(_0231_));
 sky130_fd_sc_hd__nand3_1 _0900_ (.A(_0069_),
    .B(_0231_),
    .C(net109),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _0901_ (.A(_0230_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand3_1 _0902_ (.A(_0051_),
    .B(net77),
    .C(_0071_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _0903_ (.A(_0081_),
    .B(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nor2_1 _0904_ (.A(_0233_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _0905_ (.A(_0229_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21a_1 _0906_ (.A1(net13),
    .A2(_0076_),
    .B1(_0110_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _0907_ (.A(_0237_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3_1 _0908_ (.A(_0220_),
    .B(_0239_),
    .C(_0141_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand3_1 _0909_ (.A(_0202_),
    .B(_0240_),
    .C(net262),
    .Y(_0241_));
 sky130_fd_sc_hd__nand3_1 _0910_ (.A(_0164_),
    .B(_0165_),
    .C(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand3_1 _0911_ (.A(_0060_),
    .B(_0061_),
    .C(net185),
    .Y(_0243_));
 sky130_fd_sc_hd__nand3_1 _0912_ (.A(_0170_),
    .B(_0064_),
    .C(net121),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _0913_ (.A(_0243_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand3_1 _0914_ (.A(_0094_),
    .B(_0040_),
    .C(net217),
    .Y(_0246_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(_0246_),
    .B(_0105_),
    .Y(_0247_));
 sky130_fd_sc_hd__nor2_1 _0916_ (.A(_0245_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand3_1 _0917_ (.A(_0114_),
    .B(_0054_),
    .C(net249),
    .Y(_0249_));
 sky130_fd_sc_hd__nand3_1 _0918_ (.A(_0099_),
    .B(net89),
    .C(_0118_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0919_ (.A(_0249_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand3_1 _0920_ (.A(_0036_),
    .B(net57),
    .C(_0088_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand3_1 _0921_ (.A(_0060_),
    .B(net153),
    .C(_0116_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _0922_ (.A(_0252_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _0923_ (.A(_0251_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _0924_ (.A(_0248_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__or2_1 _0925_ (.A(net25),
    .B(_0081_),
    .X(_0257_));
 sky130_fd_sc_hd__nand3_1 _0926_ (.A(_0256_),
    .B(_0138_),
    .C(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nand2_1 _0927_ (.A(_0132_),
    .B(net248),
    .Y(_0259_));
 sky130_fd_sc_hd__nand3_1 _0928_ (.A(_0170_),
    .B(_0214_),
    .C(net120),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _0929_ (.A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__o21a_1 _0930_ (.A1(net152),
    .A2(_0019_),
    .B1(_0074_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_1 _0931_ (.A(_0261_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand3_1 _0932_ (.A(_0122_),
    .B(net56),
    .C(_0118_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand3_1 _0933_ (.A(_0203_),
    .B(net88),
    .C(_0129_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3_1 _0935_ (.A(_0060_),
    .B(_0187_),
    .C(net216),
    .Y(_0267_));
 sky130_fd_sc_hd__nand3_1 _0936_ (.A(_0114_),
    .B(_0126_),
    .C(net184),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _0937_ (.A(_0267_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor2_1 _0938_ (.A(_0266_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(_0263_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21a_1 _0940_ (.A1(net24),
    .A2(_0105_),
    .B1(_0111_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _0941_ (.A(_0271_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand3_1 _0942_ (.A(_0258_),
    .B(net261),
    .C(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nand2_1 _0943_ (.A(_0132_),
    .B(net245),
    .Y(_0275_));
 sky130_fd_sc_hd__nand3_1 _0944_ (.A(_0068_),
    .B(_0051_),
    .C(net213),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_1 _0945_ (.A(_0275_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _0946_ (.A(net85),
    .Y(_0278_));
 sky130_fd_sc_hd__nand3_1 _0947_ (.A(_0094_),
    .B(_0061_),
    .C(net181),
    .Y(_0279_));
 sky130_fd_sc_hd__o21ai_1 _0948_ (.A1(_0278_),
    .A2(_0104_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _0949_ (.A(_0277_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand3_1 _0950_ (.A(_0191_),
    .B(_0057_),
    .C(net117),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0951_ (.A(_0134_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _0952_ (.A(_0074_),
    .B(net149),
    .Y(_0284_));
 sky130_fd_sc_hd__nand3_1 _0953_ (.A(_0061_),
    .B(net53),
    .C(_0064_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2_1 _0954_ (.A(_0284_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_1 _0955_ (.A(_0283_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _0956_ (.A(_0281_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21a_1 _0957_ (.A1(net21),
    .A2(_0105_),
    .B1(_0111_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _0958_ (.A(_0288_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__buf_2 _0959_ (.A(_0038_),
    .X(_0291_));
 sky130_fd_sc_hd__nand3_1 _0960_ (.A(_0068_),
    .B(_0291_),
    .C(net214),
    .Y(_0292_));
 sky130_fd_sc_hd__nand3_1 _0961_ (.A(_0191_),
    .B(_0071_),
    .C(net118),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _0962_ (.A(_0292_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand3_1 _0963_ (.A(_0098_),
    .B(_0126_),
    .C(net182),
    .Y(_0295_));
 sky130_fd_sc_hd__nand2_1 _0964_ (.A(_0295_),
    .B(_0134_),
    .Y(_0296_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(_0294_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__nand3_1 _0966_ (.A(_0222_),
    .B(_0069_),
    .C(net246),
    .Y(_0298_));
 sky130_fd_sc_hd__nand3_1 _0967_ (.A(_0093_),
    .B(net150),
    .C(_0223_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _0968_ (.A(_0298_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand3_1 _0969_ (.A(_0061_),
    .B(net54),
    .C(_0214_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand3_1 _0970_ (.A(_0203_),
    .B(net86),
    .C(_0057_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_1 _0972_ (.A(_0300_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_1 _0973_ (.A(_0297_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21a_1 _0974_ (.A1(net22),
    .A2(_0144_),
    .B1(_0138_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(_0305_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand3_1 _0976_ (.A(_0290_),
    .B(_0307_),
    .C(_0141_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand3_1 _0977_ (.A(_0274_),
    .B(net262),
    .C(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2_1 _0978_ (.A(_0132_),
    .B(net243),
    .Y(_0310_));
 sky130_fd_sc_hd__nand3_1 _0979_ (.A(_0061_),
    .B(net51),
    .C(_0214_),
    .Y(_0311_));
 sky130_fd_sc_hd__nand2_1 _0980_ (.A(_0310_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(net211),
    .Y(_0313_));
 sky130_fd_sc_hd__nand3_1 _0982_ (.A(_0094_),
    .B(net147),
    .C(_0116_),
    .Y(_0314_));
 sky130_fd_sc_hd__o21ai_1 _0983_ (.A1(_0313_),
    .A2(_0157_),
    .B1(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(_0312_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand3_1 _0985_ (.A(_0187_),
    .B(net83),
    .C(_0214_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand3_1 _0986_ (.A(_0054_),
    .B(_0127_),
    .C(net115),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(_0317_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__nand3_1 _0988_ (.A(_0060_),
    .B(_0061_),
    .C(net179),
    .Y(_0320_));
 sky130_fd_sc_hd__nand2_1 _0989_ (.A(_0320_),
    .B(_0076_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _0990_ (.A(_0319_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(_0316_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__o21a_1 _0992_ (.A1(net19),
    .A2(_0109_),
    .B1(_0111_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0323_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand3_1 _0994_ (.A(_0126_),
    .B(net52),
    .C(_0127_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand3_1 _0995_ (.A(_0222_),
    .B(net148),
    .C(_0223_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand3_1 _0997_ (.A(_0098_),
    .B(_0099_),
    .C(net212),
    .Y(_0329_));
 sky130_fd_sc_hd__nand3_1 _0998_ (.A(_0050_),
    .B(_0183_),
    .C(net180),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _0999_ (.A(_0329_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(_0328_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__buf_4 _1001_ (.A(_0049_),
    .X(_0333_));
 sky130_fd_sc_hd__nand3_1 _1002_ (.A(_0333_),
    .B(_0069_),
    .C(net244),
    .Y(_0334_));
 sky130_fd_sc_hd__nand3_1 _1003_ (.A(_0069_),
    .B(_0231_),
    .C(net116),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1004_ (.A(_0334_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand3_1 _1005_ (.A(_0203_),
    .B(net84),
    .C(_0057_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _1006_ (.A(_0134_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__nor2_1 _1007_ (.A(_0336_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(_0332_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__o21a_1 _1009_ (.A1(net20),
    .A2(_0144_),
    .B1(_0138_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _1010_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand3_1 _1011_ (.A(_0325_),
    .B(_0342_),
    .C(net261),
    .Y(_0343_));
 sky130_fd_sc_hd__nand3_1 _1012_ (.A(_0222_),
    .B(_0069_),
    .C(net241),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _1013_ (.A(_0081_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand3_1 _1014_ (.A(_0098_),
    .B(_0122_),
    .C(net177),
    .Y(_0346_));
 sky130_fd_sc_hd__nand3_1 _1015_ (.A(_0170_),
    .B(_0064_),
    .C(net113),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _1016_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nor2_1 _1017_ (.A(_0345_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand3_1 _1018_ (.A(_0051_),
    .B(net81),
    .C(_0071_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand3_1 _1019_ (.A(_0093_),
    .B(net145),
    .C(_0223_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _1020_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand3_1 _1021_ (.A(_0050_),
    .B(_0203_),
    .C(net209),
    .Y(_0353_));
 sky130_fd_sc_hd__nand3_1 _1022_ (.A(_0126_),
    .B(net49),
    .C(_0057_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _1023_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _1024_ (.A(_0352_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _1025_ (.A(_0349_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__o21a_1 _1026_ (.A1(net17),
    .A2(_0144_),
    .B1(_0110_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(_0357_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand3_1 _1028_ (.A(_0291_),
    .B(net82),
    .C(_0231_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _1029_ (.A(_0081_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand3_1 _1030_ (.A(_0068_),
    .B(_0183_),
    .C(net178),
    .Y(_0362_));
 sky130_fd_sc_hd__nand3_1 _1031_ (.A(_0333_),
    .B(_0069_),
    .C(net242),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _1033_ (.A(_0361_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand3_1 _1034_ (.A(_0093_),
    .B(net146),
    .C(_0115_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand3_1 _1035_ (.A(_0053_),
    .B(_0231_),
    .C(net114),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _1036_ (.A(_0366_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand3_1 _1037_ (.A(_0333_),
    .B(_0291_),
    .C(net210),
    .Y(_0369_));
 sky130_fd_sc_hd__nand3_1 _1038_ (.A(_0035_),
    .B(net50),
    .C(_0231_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(_0369_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _1040_ (.A(_0368_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(_0365_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__o21a_1 _1042_ (.A1(net18),
    .A2(_0134_),
    .B1(net260),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand3_1 _1044_ (.A(_0359_),
    .B(_0375_),
    .C(_0141_),
    .Y(_0376_));
 sky130_fd_sc_hd__clkinv_2 _1045_ (.A(net262),
    .Y(_0377_));
 sky130_fd_sc_hd__nand3_1 _1046_ (.A(_0343_),
    .B(_0376_),
    .C(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__nand3_1 _1047_ (.A(_0309_),
    .B(_0378_),
    .C(net263),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(_0242_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _1049_ (.A(_0380_),
    .B(net264),
    .Y(_0381_));
 sky130_fd_sc_hd__nand2_1 _1050_ (.A(_0021_),
    .B(net252),
    .Y(_0382_));
 sky130_fd_sc_hd__nand3_1 _1051_ (.A(_0040_),
    .B(net92),
    .C(_0088_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_1 _1052_ (.A(_0382_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(net188),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_2 _1054_ (.A(_0048_),
    .B(_0034_),
    .Y(_0386_));
 sky130_fd_sc_hd__clkbuf_4 _1055_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__nand3_1 _1056_ (.A(_0036_),
    .B(net60),
    .C(_0088_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_1 _1057_ (.A1(_0385_),
    .A2(_0387_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_1 _1058_ (.A(_0384_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(net124),
    .Y(_0391_));
 sky130_fd_sc_hd__nand3_1 _1060_ (.A(_0114_),
    .B(net156),
    .C(_0116_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_1 _1061_ (.A1(_0391_),
    .A2(_0092_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(net220),
    .Y(_0394_));
 sky130_fd_sc_hd__o21ai_1 _1063_ (.A1(_0394_),
    .A2(_0157_),
    .B1(_0105_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0393_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nand2_1 _1065_ (.A(_0390_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o21a_1 _1066_ (.A1(net28),
    .A2(_0109_),
    .B1(_0138_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _1067_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand3_1 _1068_ (.A(_0126_),
    .B(net59),
    .C(_0127_),
    .Y(_0400_));
 sky130_fd_sc_hd__nand2_1 _1069_ (.A(_0076_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand3_1 _1070_ (.A(_0094_),
    .B(_0040_),
    .C(net219),
    .Y(_0402_));
 sky130_fd_sc_hd__nand3_1 _1071_ (.A(_0098_),
    .B(_0122_),
    .C(net187),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _1072_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_1 _1073_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand3_1 _1074_ (.A(_0068_),
    .B(net155),
    .C(_0116_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand3_1 _1075_ (.A(_0191_),
    .B(_0129_),
    .C(net123),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _1077_ (.A(_0132_),
    .B(net251),
    .Y(_0409_));
 sky130_fd_sc_hd__nand3_1 _1078_ (.A(_0187_),
    .B(net91),
    .C(_0214_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(_0409_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__nor2_1 _1080_ (.A(_0408_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _1081_ (.A(_0405_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21a_1 _1082_ (.A1(net27),
    .A2(_0105_),
    .B1(_0111_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(_0413_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand3_1 _1084_ (.A(_0399_),
    .B(_0415_),
    .C(_0141_),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(net222),
    .Y(_0417_));
 sky130_fd_sc_hd__nand3_1 _1086_ (.A(_0040_),
    .B(net94),
    .C(_0064_),
    .Y(_0418_));
 sky130_fd_sc_hd__o21ai_1 _1087_ (.A1(_0417_),
    .A2(_0157_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(net62),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _1089_ (.A(_0021_),
    .B(net254),
    .Y(_0421_));
 sky130_fd_sc_hd__o21ai_1 _1090_ (.A1(_0420_),
    .A2(_0148_),
    .B1(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nor2_1 _1091_ (.A(_0419_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(net158),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_4 _1093_ (.A(_0049_),
    .B(_0115_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand3_1 _1094_ (.A(_0170_),
    .B(_0214_),
    .C(net126),
    .Y(_0426_));
 sky130_fd_sc_hd__o21ai_1 _1095_ (.A1(_0424_),
    .A2(_0425_),
    .B1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(net190),
    .Y(_0428_));
 sky130_fd_sc_hd__o21ai_1 _1097_ (.A1(_0428_),
    .A2(_0387_),
    .B1(_0014_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_1 _1098_ (.A(_0427_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _1099_ (.A(_0423_),
    .B(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(net221),
    .Y(_0432_));
 sky130_fd_sc_hd__nand3_1 _1101_ (.A(_0099_),
    .B(net93),
    .C(_0118_),
    .Y(_0433_));
 sky130_fd_sc_hd__o21ai_1 _1102_ (.A1(_0432_),
    .A2(_0157_),
    .B1(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(net61),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0021_),
    .B(net253),
    .Y(_0436_));
 sky130_fd_sc_hd__o21ai_1 _1105_ (.A1(_0435_),
    .A2(_0148_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(_0434_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(net157),
    .Y(_0439_));
 sky130_fd_sc_hd__nand3_1 _1108_ (.A(_0054_),
    .B(_0057_),
    .C(net125),
    .Y(_0440_));
 sky130_fd_sc_hd__o21ai_1 _1109_ (.A1(_0439_),
    .A2(_0425_),
    .B1(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _1110_ (.A(net189),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_1 _1111_ (.A1(_0442_),
    .A2(_0387_),
    .B1(_0085_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(_0441_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(_0438_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _1114_ (.A(_0431_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _1115_ (.A(_0446_),
    .B(_0109_),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_2 _1116_ (.A(_0085_),
    .Y(_0448_));
 sky130_fd_sc_hd__o22ai_1 _1117_ (.A1(net30),
    .A2(_0013_),
    .B1(net29),
    .B2(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _1118_ (.A(_0115_),
    .B(_0044_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_2 _1119_ (.A(_0450_),
    .B(_0018_),
    .Y(_0451_));
 sky130_fd_sc_hd__a21oi_1 _1120_ (.A1(_0449_),
    .A2(_0451_),
    .B1(_0377_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand3_1 _1121_ (.A(_0416_),
    .B(_0447_),
    .C(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__a21o_1 _1122_ (.A1(_0451_),
    .A2(net23),
    .B1(_0448_),
    .X(_0454_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(net151),
    .Y(_0455_));
 sky130_fd_sc_hd__nand3_1 _1124_ (.A(_0069_),
    .B(_0231_),
    .C(net119),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_1 _1125_ (.A1(_0455_),
    .A2(_0425_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(net55),
    .Y(_0458_));
 sky130_fd_sc_hd__buf_2 _1127_ (.A(_0020_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _1128_ (.A(_0459_),
    .B(net247),
    .Y(_0460_));
 sky130_fd_sc_hd__o21ai_1 _1129_ (.A1(_0458_),
    .A2(_0148_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _1130_ (.A(_0457_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand3_1 _1131_ (.A(_0039_),
    .B(net87),
    .C(_0063_),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(net183),
    .Y(_0465_));
 sky130_fd_sc_hd__nand3_1 _1134_ (.A(_0222_),
    .B(_0291_),
    .C(net215),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_1 _1135_ (.A1(_0465_),
    .A2(_0386_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__nor2_1 _1136_ (.A(_0464_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(_0462_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(_0454_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _1139_ (.A(_0459_),
    .B(net250),
    .Y(_0471_));
 sky130_fd_sc_hd__nand3_1 _1140_ (.A(_0333_),
    .B(net154),
    .C(_0223_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _1141_ (.A(_0471_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _1142_ (.A(net218),
    .Y(_0474_));
 sky130_fd_sc_hd__nand3_1 _1143_ (.A(_0170_),
    .B(_0088_),
    .C(net122),
    .Y(_0475_));
 sky130_fd_sc_hd__o21ai_1 _1144_ (.A1(_0474_),
    .A2(_0157_),
    .B1(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nor2_1 _1145_ (.A(_0473_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__and2b_1 _1146_ (.A_N(_0386_),
    .B(net186),
    .X(_0478_));
 sky130_fd_sc_hd__inv_2 _1147_ (.A(net90),
    .Y(_0479_));
 sky130_fd_sc_hd__nand3_1 _1148_ (.A(_0122_),
    .B(net58),
    .C(_0118_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_1 _1149_ (.A1(_0479_),
    .A2(_0104_),
    .B1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor2_1 _1150_ (.A(_0478_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21oi_1 _1151_ (.A1(_0451_),
    .A2(net26),
    .B1(_0013_),
    .Y(_0483_));
 sky130_fd_sc_hd__nand3_1 _1152_ (.A(_0477_),
    .B(_0482_),
    .C(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_1 _1153_ (.A(_0484_),
    .B(_0377_),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _1154_ (.A(_0470_),
    .B(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _1155_ (.A(net33),
    .Y(_0487_));
 sky130_fd_sc_hd__nand3_1 _1156_ (.A(_0170_),
    .B(_0118_),
    .C(net97),
    .Y(_0488_));
 sky130_fd_sc_hd__o21ai_1 _1157_ (.A1(_0487_),
    .A2(_0148_),
    .B1(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _1158_ (.A(net161),
    .Y(_0490_));
 sky130_fd_sc_hd__nand3_1 _1159_ (.A(_0060_),
    .B(_0099_),
    .C(net193),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_1 _1160_ (.A1(_0490_),
    .A2(_0387_),
    .B1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__nor2_1 _1161_ (.A(_0489_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _1162_ (.A(_0459_),
    .B(net225),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(_0494_),
    .B(_0081_),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(net129),
    .Y(_0496_));
 sky130_fd_sc_hd__nand3_1 _1165_ (.A(_0187_),
    .B(net65),
    .C(_0064_),
    .Y(_0497_));
 sky130_fd_sc_hd__o21ai_1 _1166_ (.A1(_0496_),
    .A2(_0425_),
    .B1(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__nor2_1 _1167_ (.A(_0495_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1168_ (.A(_0493_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21a_1 _1169_ (.A1(net1),
    .A2(_0144_),
    .B1(_0111_),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _1170_ (.A(_0500_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand3_1 _1171_ (.A(_0291_),
    .B(net76),
    .C(_0231_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(_0081_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(net172),
    .Y(_0505_));
 sky130_fd_sc_hd__nand3_1 _1174_ (.A(_0122_),
    .B(net44),
    .C(_0118_),
    .Y(_0506_));
 sky130_fd_sc_hd__o21ai_1 _1175_ (.A1(_0505_),
    .A2(_0387_),
    .B1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__nor2_1 _1176_ (.A(_0504_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(_0459_),
    .B(net236),
    .Y(_0509_));
 sky130_fd_sc_hd__nand3_1 _1178_ (.A(_0093_),
    .B(_0039_),
    .C(net204),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1179_ (.A(_0509_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(net108),
    .Y(_0512_));
 sky130_fd_sc_hd__nand3_1 _1181_ (.A(_0333_),
    .B(net140),
    .C(_0223_),
    .Y(_0513_));
 sky130_fd_sc_hd__o21ai_1 _1182_ (.A1(_0512_),
    .A2(_0092_),
    .B1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1183_ (.A(_0511_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _1184_ (.A(_0508_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__o21a_1 _1185_ (.A1(net12),
    .A2(_0076_),
    .B1(net260),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(_0516_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand3_1 _1187_ (.A(_0502_),
    .B(_0518_),
    .C(_0141_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _1188_ (.A(_0486_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand3_1 _1189_ (.A(_0453_),
    .B(_0165_),
    .C(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1190_ (.A(_0132_),
    .B(net229),
    .Y(_0522_));
 sky130_fd_sc_hd__nand3_1 _1191_ (.A(_0187_),
    .B(net69),
    .C(_0214_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(_0522_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(net165),
    .Y(_0525_));
 sky130_fd_sc_hd__nand3_1 _1194_ (.A(_0036_),
    .B(net37),
    .C(_0088_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _1195_ (.A1(_0525_),
    .A2(_0387_),
    .B1(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_1 _1196_ (.A(_0524_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand3_1 _1197_ (.A(_0050_),
    .B(net133),
    .C(_0116_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand3_1 _1198_ (.A(_0054_),
    .B(_0127_),
    .C(net101),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand3_1 _1200_ (.A(_0060_),
    .B(_0187_),
    .C(net197),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _1201_ (.A(_0532_),
    .B(_0076_),
    .Y(_0533_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(_0531_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(_0528_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21a_1 _1204_ (.A1(net5),
    .A2(_0109_),
    .B1(_0138_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand3_1 _1206_ (.A(_0183_),
    .B(net36),
    .C(_0129_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _1207_ (.A(_0134_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand3_1 _1208_ (.A(_0098_),
    .B(_0099_),
    .C(net196),
    .Y(_0540_));
 sky130_fd_sc_hd__nand3_1 _1209_ (.A(_0050_),
    .B(_0126_),
    .C(net164),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _1211_ (.A(_0539_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand3_1 _1212_ (.A(_0333_),
    .B(net132),
    .C(_0223_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand3_1 _1213_ (.A(_0191_),
    .B(_0071_),
    .C(net100),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0544_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _1215_ (.A(_0132_),
    .B(net228),
    .Y(_0547_));
 sky130_fd_sc_hd__nand3_1 _1216_ (.A(_0099_),
    .B(net68),
    .C(_0127_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _1217_ (.A(_0547_),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1218_ (.A(_0546_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2_1 _1219_ (.A(_0543_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__o21a_1 _1220_ (.A1(net4),
    .A2(_0144_),
    .B1(_0110_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _1221_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand3_1 _1222_ (.A(_0537_),
    .B(_0553_),
    .C(_0141_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _1223_ (.A(net134),
    .Y(_0555_));
 sky130_fd_sc_hd__nand3_1 _1224_ (.A(_0050_),
    .B(_0051_),
    .C(net198),
    .Y(_0556_));
 sky130_fd_sc_hd__o21ai_1 _1225_ (.A1(_0555_),
    .A2(_0425_),
    .B1(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _1226_ (.A(net38),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(_0021_),
    .B(net230),
    .Y(_0559_));
 sky130_fd_sc_hd__o21ai_1 _1228_ (.A1(_0558_),
    .A2(_0148_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__nor2_1 _1229_ (.A(_0557_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _1230_ (.A(net70),
    .Y(_0562_));
 sky130_fd_sc_hd__nand3_1 _1231_ (.A(_0054_),
    .B(_0057_),
    .C(net102),
    .Y(_0563_));
 sky130_fd_sc_hd__o21ai_1 _1232_ (.A1(_0562_),
    .A2(_0104_),
    .B1(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_2 _1233_ (.A(net166),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_1 _1234_ (.A1(_0565_),
    .A2(_0387_),
    .B1(_0085_),
    .Y(_0566_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(_0564_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(_0561_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_2 _1237_ (.A(net199),
    .Y(_0569_));
 sky130_fd_sc_hd__nand3_1 _1238_ (.A(_0203_),
    .B(net71),
    .C(_0129_),
    .Y(_0570_));
 sky130_fd_sc_hd__o21ai_1 _1239_ (.A1(_0569_),
    .A2(_0156_),
    .B1(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_2 _1240_ (.A(net39),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _1241_ (.A(_0132_),
    .B(net231),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_1 _1242_ (.A1(_0572_),
    .A2(_0148_),
    .B1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(_0571_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _1244_ (.A(net135),
    .Y(_0576_));
 sky130_fd_sc_hd__nand3_1 _1245_ (.A(_0191_),
    .B(_0071_),
    .C(net103),
    .Y(_0577_));
 sky130_fd_sc_hd__o21ai_1 _1246_ (.A1(_0576_),
    .A2(_0425_),
    .B1(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_2 _1247_ (.A(net167),
    .Y(_0579_));
 sky130_fd_sc_hd__o21ai_1 _1248_ (.A1(_0579_),
    .A2(_0386_),
    .B1(_0014_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _1249_ (.A(_0578_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(_0575_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2_1 _1251_ (.A(_0568_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0583_),
    .B(_0109_),
    .Y(_0584_));
 sky130_fd_sc_hd__o22ai_1 _1253_ (.A1(net7),
    .A2(_0013_),
    .B1(net6),
    .B2(_0448_),
    .Y(_0585_));
 sky130_fd_sc_hd__a21oi_1 _1254_ (.A1(_0585_),
    .A2(_0451_),
    .B1(_0377_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand3_1 _1255_ (.A(_0554_),
    .B(_0584_),
    .C(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__a21o_1 _1256_ (.A1(_0451_),
    .A2(net3),
    .B1(_0013_),
    .X(_0588_));
 sky130_fd_sc_hd__inv_2 _1257_ (.A(net99),
    .Y(_0589_));
 sky130_fd_sc_hd__nand3_1 _1258_ (.A(_0093_),
    .B(net131),
    .C(_0115_),
    .Y(_0590_));
 sky130_fd_sc_hd__o21ai_1 _1259_ (.A1(_0589_),
    .A2(_0092_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(net35),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _1261_ (.A(_0459_),
    .B(net227),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_1 _1262_ (.A1(_0592_),
    .A2(_0147_),
    .B1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nor2_1 _1263_ (.A(_0591_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand3_1 _1264_ (.A(_0039_),
    .B(net67),
    .C(_0056_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _1266_ (.A(net163),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3_1 _1267_ (.A(_0093_),
    .B(_0291_),
    .C(net195),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_1 _1268_ (.A1(_0598_),
    .A2(_0386_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _1269_ (.A(_0597_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_1 _1270_ (.A(_0595_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(_0588_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand3_1 _1272_ (.A(_0333_),
    .B(_0035_),
    .C(net162),
    .Y(_0604_));
 sky130_fd_sc_hd__nand3_1 _1273_ (.A(_0222_),
    .B(net130),
    .C(_0223_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(_0604_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _1275_ (.A(net194),
    .Y(_0607_));
 sky130_fd_sc_hd__nand2_1 _1276_ (.A(_0459_),
    .B(net226),
    .Y(_0608_));
 sky130_fd_sc_hd__o21ai_1 _1277_ (.A1(_0607_),
    .A2(_0157_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _1278_ (.A(_0606_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand3_1 _1279_ (.A(_0039_),
    .B(net66),
    .C(_0063_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _1280_ (.A(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _1281_ (.A(net98),
    .Y(_0613_));
 sky130_fd_sc_hd__nand3_1 _1282_ (.A(_0183_),
    .B(net34),
    .C(_0129_),
    .Y(_0614_));
 sky130_fd_sc_hd__o21ai_1 _1283_ (.A1(_0613_),
    .A2(_0092_),
    .B1(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nor2_1 _1284_ (.A(_0612_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21oi_1 _1285_ (.A1(_0451_),
    .A2(net2),
    .B1(_0448_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand3_1 _1286_ (.A(_0610_),
    .B(_0616_),
    .C(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _1287_ (.A(_0618_),
    .B(_0377_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _1288_ (.A(_0603_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__inv_2 _1289_ (.A(net63),
    .Y(_0621_));
 sky130_fd_sc_hd__nand3_1 _1290_ (.A(_0191_),
    .B(_0129_),
    .C(net127),
    .Y(_0622_));
 sky130_fd_sc_hd__o21ai_1 _1291_ (.A1(_0621_),
    .A2(_0147_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _1292_ (.A(net191),
    .Y(_0624_));
 sky130_fd_sc_hd__nand3_1 _1293_ (.A(_0114_),
    .B(_0203_),
    .C(net223),
    .Y(_0625_));
 sky130_fd_sc_hd__o21ai_1 _1294_ (.A1(_0624_),
    .A2(_0387_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nor2_1 _1295_ (.A(_0623_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(_0459_),
    .B(net255),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _1297_ (.A(_0628_),
    .B(_0081_),
    .Y(_0629_));
 sky130_fd_sc_hd__inv_2 _1298_ (.A(net159),
    .Y(_0630_));
 sky130_fd_sc_hd__nand3_1 _1299_ (.A(_0099_),
    .B(net95),
    .C(_0127_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_1 _1300_ (.A1(_0630_),
    .A2(_0425_),
    .B1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nor2_1 _1301_ (.A(_0629_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _1302_ (.A(_0627_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__o21a_1 _1303_ (.A1(net31),
    .A2(_0144_),
    .B1(_0110_),
    .X(_0635_));
 sky130_fd_sc_hd__nand2_1 _1304_ (.A(_0634_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(_0459_),
    .B(net256),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(_0637_),
    .B(_0075_),
    .Y(_0638_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(net64),
    .Y(_0639_));
 sky130_fd_sc_hd__nand3_1 _1308_ (.A(_0333_),
    .B(_0035_),
    .C(net192),
    .Y(_0640_));
 sky130_fd_sc_hd__o21ai_1 _1309_ (.A1(_0639_),
    .A2(_0148_),
    .B1(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor2_1 _1310_ (.A(_0638_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand3_1 _1311_ (.A(_0093_),
    .B(net160),
    .C(_0115_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand3_1 _1312_ (.A(_0053_),
    .B(_0063_),
    .C(net128),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _1313_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand3_1 _1314_ (.A(_0222_),
    .B(_0291_),
    .C(net224),
    .Y(_0646_));
 sky130_fd_sc_hd__nand3_1 _1315_ (.A(_0291_),
    .B(net96),
    .C(_0231_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _1316_ (.A(_0646_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__nor2_1 _1317_ (.A(_0645_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0642_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21a_1 _1319_ (.A1(net32),
    .A2(_0134_),
    .B1(net260),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _1320_ (.A(_0650_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand3_1 _1321_ (.A(_0636_),
    .B(_0652_),
    .C(_0141_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(_0620_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand3_1 _1323_ (.A(_0587_),
    .B(net263),
    .C(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(_0521_),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(net264),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _1326_ (.A(_0656_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__and3_1 _1327_ (.A(_0027_),
    .B(_0018_),
    .C(net257),
    .X(_0659_));
 sky130_fd_sc_hd__nand3_1 _1328_ (.A(_0381_),
    .B(_0658_),
    .C(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _1329_ (.A(_0028_),
    .B(net271),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _1330_ (.A(_0660_),
    .B(_0661_),
    .Y(_0005_));
 sky130_fd_sc_hd__a221o_1 _1331_ (.A1(net266),
    .A2(_0028_),
    .B1(_0016_),
    .B2(_0023_),
    .C1(_0032_),
    .X(_0006_));
 sky130_fd_sc_hd__nor2_1 _1332_ (.A(_0110_),
    .B(_0032_),
    .Y(_0662_));
 sky130_fd_sc_hd__a21oi_1 _1333_ (.A1(_0026_),
    .A2(_0111_),
    .B1(_0662_),
    .Y(_0007_));
 sky130_fd_sc_hd__a21o_1 _1334_ (.A1(_0016_),
    .A2(_0018_),
    .B1(_0025_),
    .X(_0663_));
 sky130_fd_sc_hd__inv_2 _1335_ (.A(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _1336_ (.A(_0662_),
    .B(net261),
    .Y(_0665_));
 sky130_fd_sc_hd__or2_1 _1337_ (.A(net261),
    .B(_0662_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _1338_ (.A(_0664_),
    .B(_0665_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_1 _1339_ (.A(_0667_),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_1 _1340_ (.A(_0377_),
    .B(_0665_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0665_),
    .B(_0377_),
    .Y(_0669_));
 sky130_fd_sc_hd__and3b_1 _1342_ (.A_N(_0668_),
    .B(_0664_),
    .C(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(_0670_),
    .X(_0009_));
 sky130_fd_sc_hd__nor2_1 _1344_ (.A(net263),
    .B(_0668_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0668_),
    .B(net263),
    .Y(_0672_));
 sky130_fd_sc_hd__or3b_1 _1346_ (.A(_0663_),
    .B(_0671_),
    .C_N(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(_0673_),
    .Y(_0010_));
 sky130_fd_sc_hd__a21o_1 _1348_ (.A1(_0672_),
    .A2(_0657_),
    .B1(_0663_),
    .X(_0674_));
 sky130_fd_sc_hd__inv_2 _1349_ (.A(_0674_),
    .Y(_0011_));
 sky130_fd_sc_hd__and3_1 _1350_ (.A(_0023_),
    .B(net272),
    .C(net265),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _1351_ (.A(_0675_),
    .X(_0012_));
 sky130_fd_sc_hd__dfrtp_4 _1352_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0001_),
    .RESET_B(net273),
    .Q(net267));
 sky130_fd_sc_hd__dfrtp_4 _1353_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0002_),
    .RESET_B(net273),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_4 _1354_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0003_),
    .RESET_B(net274),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_2 _1355_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0004_),
    .RESET_B(net274),
    .Q(net270));
 sky130_fd_sc_hd__dfrtp_1 _1356_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0005_),
    .RESET_B(net274),
    .Q(net271));
 sky130_fd_sc_hd__dfrtp_1 _1357_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0000_),
    .RESET_B(net274),
    .Q(net259));
 sky130_fd_sc_hd__dfrtp_1 _1358_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0006_),
    .RESET_B(net274),
    .Q(net266));
 sky130_fd_sc_hd__dfrtp_4 _1359_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0007_),
    .RESET_B(net273),
    .Q(net260));
 sky130_fd_sc_hd__dfrtp_4 _1360_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0008_),
    .RESET_B(net273),
    .Q(net261));
 sky130_fd_sc_hd__dfrtp_4 _1361_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0009_),
    .RESET_B(net273),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_4 _1362_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0010_),
    .RESET_B(net273),
    .Q(net263));
 sky130_fd_sc_hd__dfrtp_2 _1363_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0011_),
    .RESET_B(net273),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_1 _1364_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0012_),
    .RESET_B(net273),
    .Q(net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_1__leaf_CLK));
 sky130_fd_sc_hd__buf_2 fanout272 (.A(net270),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(net258),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 fanout274 (.A(net258),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(PAR_IN1[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(PAR_IN1[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(PAR_IN4[12]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(PAR_IN4[13]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(PAR_IN4[14]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(PAR_IN4[15]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(PAR_IN4[16]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(PAR_IN4[17]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(PAR_IN4[18]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(PAR_IN4[19]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(PAR_IN4[1]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(PAR_IN4[20]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(PAR_IN1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(PAR_IN4[21]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(PAR_IN4[22]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(PAR_IN4[23]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(PAR_IN4[24]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(PAR_IN4[25]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(PAR_IN4[26]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(PAR_IN4[27]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(PAR_IN4[28]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(PAR_IN4[29]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(PAR_IN4[2]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(PAR_IN1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(PAR_IN4[30]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(PAR_IN4[31]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(PAR_IN4[3]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(PAR_IN4[4]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(PAR_IN4[5]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(PAR_IN4[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(PAR_IN4[7]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(PAR_IN4[8]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(PAR_IN4[9]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(PAR_IN5[0]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(PAR_IN1[20]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(PAR_IN5[10]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(PAR_IN5[11]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(PAR_IN5[12]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(PAR_IN5[13]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(PAR_IN5[14]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(PAR_IN5[15]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(PAR_IN5[16]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(PAR_IN5[17]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(PAR_IN5[18]),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 input139 (.A(PAR_IN5[19]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(PAR_IN1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(PAR_IN5[1]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(PAR_IN5[20]),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 input142 (.A(PAR_IN5[21]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(PAR_IN5[22]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(PAR_IN5[23]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(PAR_IN5[24]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(PAR_IN5[25]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(PAR_IN5[26]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(PAR_IN5[27]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(PAR_IN5[28]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(PAR_IN1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(PAR_IN5[29]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(PAR_IN5[2]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(PAR_IN5[30]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(PAR_IN5[31]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(PAR_IN5[3]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(PAR_IN5[4]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(PAR_IN5[5]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(PAR_IN5[6]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(PAR_IN5[7]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(PAR_IN5[8]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(PAR_IN1[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(PAR_IN5[9]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(PAR_IN6[0]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(PAR_IN6[10]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(PAR_IN6[11]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(PAR_IN6[12]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(PAR_IN6[13]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(PAR_IN6[14]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(PAR_IN6[15]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(PAR_IN6[16]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(PAR_IN6[17]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(PAR_IN1[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(PAR_IN6[18]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(PAR_IN6[19]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(PAR_IN6[1]),
    .X(net172));
 sky130_fd_sc_hd__dlymetal6s2s_1 input173 (.A(PAR_IN6[20]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(PAR_IN6[21]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(PAR_IN6[22]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(PAR_IN6[23]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(PAR_IN6[24]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(PAR_IN6[25]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(PAR_IN6[26]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(PAR_IN1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(PAR_IN6[27]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(PAR_IN6[28]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(PAR_IN6[29]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(PAR_IN6[2]),
    .X(net183));
 sky130_fd_sc_hd__dlymetal6s2s_1 input184 (.A(PAR_IN6[30]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(PAR_IN6[31]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(PAR_IN6[3]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(PAR_IN6[4]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(PAR_IN6[5]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(PAR_IN6[6]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(PAR_IN1[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(PAR_IN6[7]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(PAR_IN6[8]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(PAR_IN6[9]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(PAR_IN7[0]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(PAR_IN7[10]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(PAR_IN7[11]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(PAR_IN7[12]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(PAR_IN7[13]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(PAR_IN7[14]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(PAR_IN7[15]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(PAR_IN1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(PAR_IN1[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(PAR_IN7[16]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(PAR_IN7[17]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(PAR_IN7[18]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(PAR_IN7[19]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(PAR_IN7[1]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(PAR_IN7[20]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(PAR_IN7[21]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(PAR_IN7[22]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(PAR_IN7[23]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(PAR_IN7[24]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(PAR_IN1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(PAR_IN7[25]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(PAR_IN7[26]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(PAR_IN7[27]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(PAR_IN7[28]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(PAR_IN7[29]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(PAR_IN7[2]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(PAR_IN7[30]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(PAR_IN7[31]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(PAR_IN7[3]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(PAR_IN7[4]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(PAR_IN1[29]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input220 (.A(PAR_IN7[5]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(PAR_IN7[6]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(PAR_IN7[7]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(PAR_IN7[8]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(PAR_IN7[9]),
    .X(net224));
 sky130_fd_sc_hd__dlymetal6s2s_1 input225 (.A(PAR_IN8[0]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(PAR_IN8[10]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(PAR_IN8[11]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(PAR_IN8[12]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(PAR_IN8[13]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(PAR_IN1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(PAR_IN8[14]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(PAR_IN8[15]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(PAR_IN8[16]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(PAR_IN8[17]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(PAR_IN8[18]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(PAR_IN8[19]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(PAR_IN8[1]),
    .X(net236));
 sky130_fd_sc_hd__dlymetal6s2s_1 input237 (.A(PAR_IN8[20]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(PAR_IN8[21]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(PAR_IN8[22]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(PAR_IN1[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(PAR_IN8[23]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(PAR_IN8[24]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(PAR_IN8[25]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(PAR_IN8[26]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(PAR_IN8[27]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 input245 (.A(PAR_IN8[28]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(PAR_IN8[29]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 input247 (.A(PAR_IN8[2]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(PAR_IN8[30]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(PAR_IN8[31]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(PAR_IN1[31]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input250 (.A(PAR_IN8[3]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(PAR_IN8[4]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(PAR_IN8[5]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(PAR_IN8[6]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(PAR_IN8[7]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(PAR_IN8[8]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(PAR_IN8[9]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 input257 (.A(READY),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 input258 (.A(RESET),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(PAR_IN1[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(PAR_IN1[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(PAR_IN1[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(PAR_IN1[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(PAR_IN1[11]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(PAR_IN1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(PAR_IN1[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(PAR_IN1[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(PAR_IN2[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(PAR_IN2[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(PAR_IN2[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(PAR_IN2[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(PAR_IN2[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(PAR_IN2[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(PAR_IN2[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(PAR_IN1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(PAR_IN2[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(PAR_IN2[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(PAR_IN2[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(PAR_IN2[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(PAR_IN2[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(PAR_IN2[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(PAR_IN2[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(PAR_IN2[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(PAR_IN2[23]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(PAR_IN2[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(PAR_IN1[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(PAR_IN2[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(PAR_IN2[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(PAR_IN2[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(PAR_IN2[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(PAR_IN2[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(PAR_IN2[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(PAR_IN2[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(PAR_IN2[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(PAR_IN2[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(PAR_IN2[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(PAR_IN1[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(PAR_IN2[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(PAR_IN2[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(PAR_IN2[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(PAR_IN2[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(PAR_IN2[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(PAR_IN3[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(PAR_IN3[10]),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 input67 (.A(PAR_IN3[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(PAR_IN3[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(PAR_IN3[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(PAR_IN1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(PAR_IN3[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(PAR_IN3[15]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(PAR_IN3[16]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(PAR_IN3[17]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(PAR_IN3[18]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(PAR_IN3[19]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(PAR_IN3[1]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(PAR_IN3[20]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(PAR_IN3[21]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(PAR_IN3[22]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(PAR_IN1[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(PAR_IN3[23]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(PAR_IN3[24]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(PAR_IN3[25]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(PAR_IN3[26]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(PAR_IN3[27]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(PAR_IN3[28]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(PAR_IN3[29]),
    .X(net86));
 sky130_fd_sc_hd__dlymetal6s2s_1 input87 (.A(PAR_IN3[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(PAR_IN3[30]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(PAR_IN3[31]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(PAR_IN1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(PAR_IN3[3]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(PAR_IN3[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(PAR_IN3[5]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(PAR_IN3[6]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(PAR_IN3[7]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(PAR_IN3[8]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(PAR_IN3[9]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(PAR_IN4[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(PAR_IN4[10]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(PAR_IN4[11]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(COMPLETE));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(COUNT[0]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(COUNT[1]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(COUNT[2]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(COUNT[3]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(COUNT[4]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(COUNT[5]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(INTERNAL_FINISH));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(SAMPLE_COUNT[0]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(SAMPLE_COUNT[1]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(SAMPLE_COUNT[2]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(SAMPLE_COUNT[3]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(SERIAL_OUT));
endmodule

