../../../../designs/lp_tree_serializer/src/lp_tree_serializer_final.sv