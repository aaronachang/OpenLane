../conv_tree_serializer/src/conv_tree_serializer.v