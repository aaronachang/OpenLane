../conv_tree_serializer/src/conv_serializer.v