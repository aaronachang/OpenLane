// This is the unpowered netlist.
module conv_tree_serializer (CLK,
    RESET,
    SERIAL_OUT,
    PAR_IN);
 input CLK;
 input RESET;
 output SERIAL_OUT;
 input [255:0] PAR_IN;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1290_;
 wire _1291_;
 wire _1294_;
 wire _1295_;
 wire _1301_;
 wire _1302_;
 wire _1305_;
 wire _1312_;
 wire _1313_;
 wire _1316_;
 wire _1323_;
 wire _1324_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1345_;
 wire _1346_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire clknet_0_CLK;
 wire clknet_0__1286_;
 wire clknet_0__1290_;
 wire clknet_0__2017_;
 wire clknet_0__2018_;
 wire clknet_0__2022_;
 wire clknet_0__2023_;
 wire clknet_0__2236_;
 wire clknet_0__2678_;
 wire clknet_0__2681_;
 wire clknet_0__2683_;
 wire clknet_0__2684_;
 wire clknet_0__2695_;
 wire clknet_0__2703_;
 wire clknet_0__2706_;
 wire clknet_0__2721_;
 wire clknet_0__2724_;
 wire clknet_0__2727_;
 wire clknet_0__2730_;
 wire clknet_0__2763_;
 wire clknet_0__2766_;
 wire clknet_0__2768_;
 wire clknet_0__2800_;
 wire clknet_0__2803_;
 wire clknet_0__2805_;
 wire clknet_0__2830_;
 wire clknet_0__2858_;
 wire clknet_1_0__leaf__1286_;
 wire clknet_1_0__leaf__1290_;
 wire clknet_1_0__leaf__2017_;
 wire clknet_1_0__leaf__2018_;
 wire clknet_1_0__leaf__2022_;
 wire clknet_1_0__leaf__2023_;
 wire clknet_1_0__leaf__2236_;
 wire clknet_1_0__leaf__2678_;
 wire clknet_1_0__leaf__2681_;
 wire clknet_1_0__leaf__2683_;
 wire clknet_1_0__leaf__2684_;
 wire clknet_1_0__leaf__2695_;
 wire clknet_1_0__leaf__2703_;
 wire clknet_1_0__leaf__2706_;
 wire clknet_1_0__leaf__2721_;
 wire clknet_1_0__leaf__2724_;
 wire clknet_1_0__leaf__2727_;
 wire clknet_1_0__leaf__2730_;
 wire clknet_1_0__leaf__2763_;
 wire clknet_1_0__leaf__2766_;
 wire clknet_1_0__leaf__2768_;
 wire clknet_1_0__leaf__2800_;
 wire clknet_1_0__leaf__2803_;
 wire clknet_1_0__leaf__2805_;
 wire clknet_1_0__leaf__2830_;
 wire clknet_1_0__leaf__2858_;
 wire clknet_1_1__leaf__1286_;
 wire clknet_1_1__leaf__1290_;
 wire clknet_1_1__leaf__2017_;
 wire clknet_1_1__leaf__2018_;
 wire clknet_1_1__leaf__2022_;
 wire clknet_1_1__leaf__2023_;
 wire clknet_1_1__leaf__2236_;
 wire clknet_1_1__leaf__2678_;
 wire clknet_1_1__leaf__2681_;
 wire clknet_1_1__leaf__2683_;
 wire clknet_1_1__leaf__2684_;
 wire clknet_1_1__leaf__2695_;
 wire clknet_1_1__leaf__2703_;
 wire clknet_1_1__leaf__2706_;
 wire clknet_1_1__leaf__2721_;
 wire clknet_1_1__leaf__2724_;
 wire clknet_1_1__leaf__2727_;
 wire clknet_1_1__leaf__2730_;
 wire clknet_1_1__leaf__2763_;
 wire clknet_1_1__leaf__2766_;
 wire clknet_1_1__leaf__2768_;
 wire clknet_1_1__leaf__2800_;
 wire clknet_1_1__leaf__2803_;
 wire clknet_1_1__leaf__2805_;
 wire clknet_1_1__leaf__2830_;
 wire clknet_1_1__leaf__2858_;
 wire clknet_3_0__leaf_CLK;
 wire clknet_3_1__leaf_CLK;
 wire clknet_3_2__leaf_CLK;
 wire clknet_3_3__leaf_CLK;
 wire clknet_3_4__leaf_CLK;
 wire clknet_3_5__leaf_CLK;
 wire clknet_3_6__leaf_CLK;
 wire clknet_3_7__leaf_CLK;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \stage_gen[1].genblk1.clks.clk_o ;
 wire \stage_gen[1].genblk1.clks.counter[0] ;
 wire \stage_gen[1].genblk1.clks.counter[1] ;
 wire \stage_gen[1].genblk1.clks.counter[2] ;
 wire \stage_gen[1].genblk1.clks.counter[3] ;
 wire \stage_gen[1].genblk1.clks.counter[4] ;
 wire \stage_gen[1].genblk1.clks.counter[5] ;
 wire \stage_gen[1].genblk1.clks.counter[6] ;
 wire \stage_gen[1].genblk1.clks.counter[7] ;
 wire \stage_gen[1].genblk1.clks.counter[8] ;
 wire \stage_gen[1].genblk1.clks.counter[9] ;
 wire \stage_gen[1].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[100].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[100].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[100].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[100].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[100].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[101].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[101].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[101].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[101].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[101].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[102].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[102].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[102].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[102].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[102].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[103].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[103].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[103].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[103].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[103].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[104].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[104].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[104].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[104].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[104].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[105].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[105].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[105].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[105].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[105].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[106].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[106].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[106].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[106].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[106].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[107].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[107].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[107].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[107].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[107].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[108].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[108].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[108].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[108].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[108].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[109].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[109].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[109].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[109].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[109].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[10].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[10].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[10].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[10].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[10].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[110].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[110].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[110].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[110].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[110].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[111].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[111].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[111].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[111].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[111].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[112].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[112].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[112].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[112].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[112].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[113].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[113].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[113].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[113].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[113].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[114].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[114].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[114].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[114].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[114].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[115].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[115].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[115].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[115].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[115].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[116].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[116].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[116].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[116].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[116].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[117].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[117].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[117].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[117].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[117].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[118].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[118].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[118].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[118].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[118].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[119].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[119].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[119].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[119].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[119].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[11].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[11].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[11].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[11].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[11].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[120].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[120].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[120].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[120].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[120].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[121].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[121].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[121].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[121].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[121].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[122].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[122].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[122].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[122].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[122].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[123].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[123].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[123].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[123].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[123].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[124].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[124].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[124].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[124].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[124].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[125].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[125].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[125].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[125].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[125].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[126].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[126].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[126].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[126].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[126].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[127].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[127].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[127].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[127].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[127].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[12].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[12].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[12].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[12].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[12].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[13].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[13].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[13].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[13].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[13].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[14].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[14].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[14].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[14].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[14].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[15].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[15].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[15].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[15].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[15].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[16].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[16].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[16].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[16].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[16].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[17].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[17].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[17].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[17].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[17].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[18].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[18].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[18].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[18].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[18].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[19].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[19].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[19].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[19].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[19].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[20].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[20].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[20].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[20].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[20].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[21].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[21].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[21].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[21].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[21].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[22].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[22].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[22].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[22].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[22].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[23].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[23].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[23].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[23].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[23].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[24].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[24].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[24].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[24].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[24].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[25].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[25].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[25].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[25].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[25].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[26].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[26].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[26].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[26].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[26].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[27].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[27].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[27].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[27].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[27].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[28].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[28].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[28].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[28].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[28].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[29].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[29].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[29].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[29].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[29].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[30].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[30].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[30].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[30].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[30].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[31].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[31].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[31].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[31].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[31].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[32].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[32].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[32].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[32].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[32].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[33].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[33].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[33].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[33].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[33].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[34].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[34].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[34].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[34].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[34].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[35].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[35].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[35].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[35].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[35].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[36].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[36].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[36].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[36].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[36].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[37].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[37].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[37].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[37].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[37].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[38].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[38].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[38].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[38].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[38].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[39].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[39].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[39].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[39].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[39].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[40].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[40].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[40].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[40].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[40].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[41].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[41].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[41].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[41].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[41].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[42].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[42].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[42].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[42].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[42].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[43].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[43].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[43].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[43].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[43].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[44].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[44].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[44].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[44].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[44].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[45].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[45].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[45].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[45].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[45].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[46].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[46].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[46].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[46].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[46].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[47].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[47].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[47].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[47].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[47].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[48].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[48].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[48].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[48].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[48].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[49].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[49].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[49].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[49].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[49].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[4].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[4].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[4].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[4].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[4].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[50].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[50].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[50].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[50].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[50].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[51].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[51].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[51].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[51].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[51].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[52].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[52].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[52].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[52].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[52].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[53].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[53].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[53].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[53].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[53].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[54].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[54].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[54].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[54].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[54].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[55].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[55].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[55].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[55].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[55].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[56].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[56].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[56].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[56].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[56].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[57].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[57].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[57].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[57].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[57].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[58].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[58].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[58].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[58].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[58].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[59].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[59].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[59].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[59].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[59].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[5].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[5].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[5].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[5].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[5].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[60].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[60].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[60].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[60].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[60].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[61].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[61].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[61].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[61].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[61].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[62].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[62].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[62].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[62].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[62].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[63].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[63].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[63].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[63].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[63].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[64].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[64].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[64].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[64].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[64].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[65].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[65].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[65].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[65].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[65].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[66].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[66].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[66].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[66].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[66].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[67].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[67].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[67].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[67].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[67].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[68].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[68].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[68].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[68].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[68].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[69].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[69].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[69].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[69].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[69].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[6].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[6].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[6].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[6].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[6].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[70].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[70].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[70].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[70].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[70].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[71].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[71].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[71].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[71].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[71].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[72].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[72].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[72].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[72].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[72].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[73].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[73].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[73].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[73].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[73].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[74].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[74].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[74].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[74].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[74].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[75].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[75].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[75].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[75].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[75].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[76].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[76].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[76].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[76].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[76].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[77].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[77].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[77].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[77].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[77].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[78].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[78].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[78].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[78].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[78].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[79].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[79].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[79].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[79].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[79].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[7].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[7].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[7].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[7].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[7].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[80].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[80].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[80].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[80].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[80].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[81].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[81].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[81].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[81].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[81].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[82].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[82].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[82].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[82].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[82].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[83].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[83].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[83].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[83].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[83].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[84].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[84].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[84].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[84].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[84].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[85].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[85].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[85].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[85].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[85].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[86].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[86].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[86].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[86].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[86].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[87].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[87].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[87].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[87].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[87].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[88].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[88].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[88].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[88].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[88].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[89].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[89].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[89].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[89].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[89].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[8].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[8].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[8].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[8].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[8].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[90].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[90].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[90].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[90].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[90].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[91].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[91].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[91].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[91].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[91].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[92].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[92].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[92].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[92].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[92].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[93].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[93].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[93].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[93].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[93].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[94].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[94].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[94].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[94].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[94].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[95].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[95].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[95].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[95].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[95].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[96].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[96].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[96].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[96].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[96].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[97].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[97].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[97].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[97].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[97].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[98].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[98].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[98].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[98].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[98].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[99].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[99].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[99].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[99].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[99].S.IN1_L5 ;
 wire \stage_gen[1].mux_gen[9].S.IN1_L1 ;
 wire \stage_gen[1].mux_gen[9].S.IN1_L2 ;
 wire \stage_gen[1].mux_gen[9].S.IN1_L3 ;
 wire \stage_gen[1].mux_gen[9].S.IN1_L4 ;
 wire \stage_gen[1].mux_gen[9].S.IN1_L5 ;
 wire \stage_gen[2].genblk1.clks.clk_o ;
 wire \stage_gen[2].genblk1.clks.counter[0] ;
 wire \stage_gen[2].genblk1.clks.counter[1] ;
 wire \stage_gen[2].genblk1.clks.counter[2] ;
 wire \stage_gen[2].genblk1.clks.counter[3] ;
 wire \stage_gen[2].genblk1.clks.counter[4] ;
 wire \stage_gen[2].genblk1.clks.counter[5] ;
 wire \stage_gen[2].genblk1.clks.counter[6] ;
 wire \stage_gen[2].genblk1.clks.counter[7] ;
 wire \stage_gen[2].genblk1.clks.counter[8] ;
 wire \stage_gen[2].genblk1.clks.counter[9] ;
 wire \stage_gen[2].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[10].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[10].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[10].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[10].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[10].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[11].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[11].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[11].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[11].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[11].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[12].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[12].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[12].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[12].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[12].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[13].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[13].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[13].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[13].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[13].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[14].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[14].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[14].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[14].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[14].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[15].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[15].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[15].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[15].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[15].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[16].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[16].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[16].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[16].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[16].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[17].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[17].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[17].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[17].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[17].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[18].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[18].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[18].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[18].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[18].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[19].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[19].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[19].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[19].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[19].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[20].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[20].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[20].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[20].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[20].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[21].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[21].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[21].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[21].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[21].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[22].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[22].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[22].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[22].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[22].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[23].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[23].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[23].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[23].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[23].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[24].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[24].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[24].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[24].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[24].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[25].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[25].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[25].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[25].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[25].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[26].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[26].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[26].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[26].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[26].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[27].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[27].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[27].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[27].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[27].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[28].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[28].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[28].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[28].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[28].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[29].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[29].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[29].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[29].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[29].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[30].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[30].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[30].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[30].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[30].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[31].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[31].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[31].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[31].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[31].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[32].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[32].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[32].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[32].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[32].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[33].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[33].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[33].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[33].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[33].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[34].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[34].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[34].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[34].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[34].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[35].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[35].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[35].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[35].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[35].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[36].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[36].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[36].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[36].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[36].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[37].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[37].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[37].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[37].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[37].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[38].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[38].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[38].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[38].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[38].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[39].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[39].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[39].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[39].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[39].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[40].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[40].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[40].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[40].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[40].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[41].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[41].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[41].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[41].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[41].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[42].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[42].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[42].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[42].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[42].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[43].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[43].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[43].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[43].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[43].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[44].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[44].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[44].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[44].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[44].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[45].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[45].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[45].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[45].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[45].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[46].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[46].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[46].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[46].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[46].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[47].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[47].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[47].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[47].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[47].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[48].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[48].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[48].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[48].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[48].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[49].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[49].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[49].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[49].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[49].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[4].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[4].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[4].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[4].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[4].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[50].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[50].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[50].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[50].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[50].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[51].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[51].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[51].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[51].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[51].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[52].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[52].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[52].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[52].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[52].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[53].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[53].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[53].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[53].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[53].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[54].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[54].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[54].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[54].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[54].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[55].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[55].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[55].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[55].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[55].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[56].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[56].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[56].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[56].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[56].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[57].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[57].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[57].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[57].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[57].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[58].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[58].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[58].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[58].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[58].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[59].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[59].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[59].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[59].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[59].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[5].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[5].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[5].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[5].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[5].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[60].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[60].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[60].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[60].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[60].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[61].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[61].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[61].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[61].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[61].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[62].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[62].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[62].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[62].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[62].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[63].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[63].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[63].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[63].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[63].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[6].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[6].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[6].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[6].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[6].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[7].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[7].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[7].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[7].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[7].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[8].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[8].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[8].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[8].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[8].S.IN1_L5 ;
 wire \stage_gen[2].mux_gen[9].S.IN1_L1 ;
 wire \stage_gen[2].mux_gen[9].S.IN1_L2 ;
 wire \stage_gen[2].mux_gen[9].S.IN1_L3 ;
 wire \stage_gen[2].mux_gen[9].S.IN1_L4 ;
 wire \stage_gen[2].mux_gen[9].S.IN1_L5 ;
 wire \stage_gen[3].genblk1.clks.clk_o ;
 wire \stage_gen[3].genblk1.clks.counter[0] ;
 wire \stage_gen[3].genblk1.clks.counter[1] ;
 wire \stage_gen[3].genblk1.clks.counter[2] ;
 wire \stage_gen[3].genblk1.clks.counter[3] ;
 wire \stage_gen[3].genblk1.clks.counter[4] ;
 wire \stage_gen[3].genblk1.clks.counter[5] ;
 wire \stage_gen[3].genblk1.clks.counter[6] ;
 wire \stage_gen[3].genblk1.clks.counter[7] ;
 wire \stage_gen[3].genblk1.clks.counter[8] ;
 wire \stage_gen[3].genblk1.clks.counter[9] ;
 wire \stage_gen[3].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[10].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[10].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[10].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[10].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[10].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[11].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[11].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[11].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[11].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[11].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[12].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[12].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[12].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[12].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[12].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[13].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[13].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[13].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[13].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[13].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[14].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[14].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[14].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[14].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[14].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[15].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[15].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[15].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[15].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[15].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[16].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[16].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[16].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[16].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[16].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[17].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[17].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[17].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[17].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[17].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[18].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[18].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[18].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[18].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[18].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[19].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[19].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[19].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[19].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[19].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[20].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[20].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[20].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[20].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[20].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[21].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[21].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[21].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[21].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[21].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[22].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[22].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[22].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[22].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[22].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[23].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[23].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[23].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[23].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[23].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[24].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[24].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[24].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[24].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[24].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[25].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[25].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[25].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[25].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[25].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[26].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[26].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[26].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[26].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[26].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[27].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[27].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[27].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[27].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[27].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[28].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[28].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[28].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[28].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[28].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[29].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[29].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[29].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[29].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[29].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[30].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[30].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[30].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[30].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[30].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[31].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[31].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[31].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[31].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[31].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[4].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[4].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[4].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[4].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[4].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[5].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[5].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[5].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[5].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[5].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[6].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[6].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[6].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[6].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[6].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[7].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[7].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[7].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[7].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[7].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[8].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[8].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[8].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[8].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[8].S.IN1_L5 ;
 wire \stage_gen[3].mux_gen[9].S.IN1_L1 ;
 wire \stage_gen[3].mux_gen[9].S.IN1_L2 ;
 wire \stage_gen[3].mux_gen[9].S.IN1_L3 ;
 wire \stage_gen[3].mux_gen[9].S.IN1_L4 ;
 wire \stage_gen[3].mux_gen[9].S.IN1_L5 ;
 wire \stage_gen[4].genblk1.clks.clk_o ;
 wire \stage_gen[4].genblk1.clks.counter[0] ;
 wire \stage_gen[4].genblk1.clks.counter[1] ;
 wire \stage_gen[4].genblk1.clks.counter[2] ;
 wire \stage_gen[4].genblk1.clks.counter[3] ;
 wire \stage_gen[4].genblk1.clks.counter[4] ;
 wire \stage_gen[4].genblk1.clks.counter[5] ;
 wire \stage_gen[4].genblk1.clks.counter[6] ;
 wire \stage_gen[4].genblk1.clks.counter[7] ;
 wire \stage_gen[4].genblk1.clks.counter[8] ;
 wire \stage_gen[4].genblk1.clks.counter[9] ;
 wire \stage_gen[4].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[10].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[10].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[10].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[10].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[10].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[11].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[11].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[11].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[11].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[11].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[12].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[12].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[12].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[12].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[12].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[13].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[13].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[13].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[13].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[13].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[14].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[14].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[14].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[14].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[14].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[15].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[15].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[15].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[15].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[15].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[4].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[4].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[4].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[4].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[4].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[5].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[5].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[5].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[5].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[5].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[6].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[6].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[6].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[6].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[6].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[7].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[7].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[7].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[7].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[7].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[8].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[8].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[8].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[8].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[8].S.IN1_L5 ;
 wire \stage_gen[4].mux_gen[9].S.IN1_L1 ;
 wire \stage_gen[4].mux_gen[9].S.IN1_L2 ;
 wire \stage_gen[4].mux_gen[9].S.IN1_L3 ;
 wire \stage_gen[4].mux_gen[9].S.IN1_L4 ;
 wire \stage_gen[4].mux_gen[9].S.IN1_L5 ;
 wire \stage_gen[5].genblk1.clks.clk_o ;
 wire \stage_gen[5].genblk1.clks.counter[0] ;
 wire \stage_gen[5].genblk1.clks.counter[1] ;
 wire \stage_gen[5].genblk1.clks.counter[2] ;
 wire \stage_gen[5].genblk1.clks.counter[3] ;
 wire \stage_gen[5].genblk1.clks.counter[4] ;
 wire \stage_gen[5].genblk1.clks.counter[5] ;
 wire \stage_gen[5].genblk1.clks.counter[6] ;
 wire \stage_gen[5].genblk1.clks.counter[7] ;
 wire \stage_gen[5].genblk1.clks.counter[8] ;
 wire \stage_gen[5].genblk1.clks.counter[9] ;
 wire \stage_gen[5].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[4].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[4].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[4].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[4].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[4].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[5].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[5].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[5].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[5].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[5].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[6].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[6].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[6].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[6].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[6].S.IN1_L5 ;
 wire \stage_gen[5].mux_gen[7].S.IN1_L1 ;
 wire \stage_gen[5].mux_gen[7].S.IN1_L2 ;
 wire \stage_gen[5].mux_gen[7].S.IN1_L3 ;
 wire \stage_gen[5].mux_gen[7].S.IN1_L4 ;
 wire \stage_gen[5].mux_gen[7].S.IN1_L5 ;
 wire \stage_gen[6].genblk1.clks.clk_o ;
 wire \stage_gen[6].genblk1.clks.counter[0] ;
 wire \stage_gen[6].genblk1.clks.counter[1] ;
 wire \stage_gen[6].genblk1.clks.counter[2] ;
 wire \stage_gen[6].genblk1.clks.counter[3] ;
 wire \stage_gen[6].genblk1.clks.counter[4] ;
 wire \stage_gen[6].genblk1.clks.counter[5] ;
 wire \stage_gen[6].genblk1.clks.counter[6] ;
 wire \stage_gen[6].genblk1.clks.counter[7] ;
 wire \stage_gen[6].genblk1.clks.counter[8] ;
 wire \stage_gen[6].genblk1.clks.counter[9] ;
 wire \stage_gen[6].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[6].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[6].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[6].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[6].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[6].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[6].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[6].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[6].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[6].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[6].mux_gen[2].S.IN1_L1 ;
 wire \stage_gen[6].mux_gen[2].S.IN1_L2 ;
 wire \stage_gen[6].mux_gen[2].S.IN1_L3 ;
 wire \stage_gen[6].mux_gen[2].S.IN1_L4 ;
 wire \stage_gen[6].mux_gen[2].S.IN1_L5 ;
 wire \stage_gen[6].mux_gen[3].S.IN1_L1 ;
 wire \stage_gen[6].mux_gen[3].S.IN1_L2 ;
 wire \stage_gen[6].mux_gen[3].S.IN1_L3 ;
 wire \stage_gen[6].mux_gen[3].S.IN1_L4 ;
 wire \stage_gen[6].mux_gen[3].S.IN1_L5 ;
 wire \stage_gen[7].genblk1.clks.clk_o ;
 wire \stage_gen[7].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[7].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[7].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[7].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[7].mux_gen[0].S.IN1_L5 ;
 wire \stage_gen[7].mux_gen[1].S.IN1_L1 ;
 wire \stage_gen[7].mux_gen[1].S.IN1_L2 ;
 wire \stage_gen[7].mux_gen[1].S.IN1_L3 ;
 wire \stage_gen[7].mux_gen[1].S.IN1_L4 ;
 wire \stage_gen[7].mux_gen[1].S.IN1_L5 ;
 wire \stage_gen[8].mux_gen[0].S.IN1_L1 ;
 wire \stage_gen[8].mux_gen[0].S.IN1_L2 ;
 wire \stage_gen[8].mux_gen[0].S.IN1_L3 ;
 wire \stage_gen[8].mux_gen[0].S.IN1_L4 ;
 wire \stage_gen[8].mux_gen[0].S.IN1_L5 ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(PAR_IN[210]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_2753_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(PAR_IN[222]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_2164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2714_));
 sky130_fd_sc_hd__decap_8 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2872_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .Y(_1358_));
 sky130_fd_sc_hd__clkbuf_4 _2873_ (.A(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__buf_6 _2874_ (.A(net257),
    .X(_1360_));
 sky130_fd_sc_hd__buf_8 _2875_ (.A(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__and3_1 _2876_ (.A(_1359_),
    .B(\stage_gen[2].mux_gen[38].S.IN1_L2 ),
    .C(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1362_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_4 _2878_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_2 _2879_ (.A(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__buf_4 _2880_ (.A(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__buf_4 _2881_ (.A(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nand2_1 _2882_ (.A(\stage_gen[1].genblk1.clks.clk_o ),
    .B(net257),
    .Y(_1367_));
 sky130_fd_sc_hd__clkinv_2 _2883_ (.A(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__buf_4 _2884_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__buf_6 _2885_ (.A(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__inv_2 _2886_ (.A(\stage_gen[1].genblk1.clks.clk_o ),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _2887_ (.A(_1371_),
    .B(net257),
    .Y(_1372_));
 sky130_fd_sc_hd__clkinv_2 _2888_ (.A(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__clkbuf_8 _2889_ (.A(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__buf_6 _2890_ (.A(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__a22oi_1 _2891_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[77].S.IN1_L5 ),
    .B1(_1375_),
    .B2(\stage_gen[1].mux_gen[77].S.IN1_L3 ),
    .Y(_1376_));
 sky130_fd_sc_hd__buf_6 _2892_ (.A(_1360_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_2 _2893_ (.A(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__and3_1 _2894_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[38].S.IN1_L4 ),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_1379_),
    .X(_0803_));
 sky130_fd_sc_hd__o21bai_1 _2896_ (.A1(_1366_),
    .A2(_1376_),
    .B1_N(_0803_),
    .Y(_0802_));
 sky130_fd_sc_hd__clkbuf_4 _2897_ (.A(_1364_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_4 _2898_ (.A(_1369_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_4 _2899_ (.A(_1374_),
    .X(_1382_));
 sky130_fd_sc_hd__a22oi_1 _2900_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[78].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[78].S.IN1_L3 ),
    .Y(_1383_));
 sky130_fd_sc_hd__buf_6 _2901_ (.A(net257),
    .X(_1384_));
 sky130_fd_sc_hd__nand2_1 _2902_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__inv_2 _2903_ (.A(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__buf_6 _2904_ (.A(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__buf_4 _2905_ (.A(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__nand2_1 _2906_ (.A(_1388_),
    .B(\stage_gen[2].mux_gen[39].S.IN1_L1 ),
    .Y(_1389_));
 sky130_fd_sc_hd__o21ai_1 _2907_ (.A1(_1380_),
    .A2(_1383_),
    .B1(_1389_),
    .Y(_0804_));
 sky130_fd_sc_hd__clkbuf_2 _2908_ (.A(net257),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _2909_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[39].S.IN1_L2 ),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1391_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2b_1 _2911_ (.A_N(_0806_),
    .B(_1389_),
    .Y(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1392_),
    .X(_0805_));
 sky130_fd_sc_hd__a22oi_1 _2913_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[79].S.IN1_L5 ),
    .B1(_1375_),
    .B2(\stage_gen[1].mux_gen[79].S.IN1_L3 ),
    .Y(_1393_));
 sky130_fd_sc_hd__and3_1 _2914_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[39].S.IN1_L4 ),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _2915_ (.A(_1394_),
    .X(_0808_));
 sky130_fd_sc_hd__o21bai_1 _2916_ (.A1(_1366_),
    .A2(_1393_),
    .B1_N(_0808_),
    .Y(_0807_));
 sky130_fd_sc_hd__a22oi_1 _2917_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[80].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[80].S.IN1_L3 ),
    .Y(_1395_));
 sky130_fd_sc_hd__nand2_1 _2918_ (.A(_1388_),
    .B(\stage_gen[2].mux_gen[40].S.IN1_L1 ),
    .Y(_1396_));
 sky130_fd_sc_hd__o21ai_1 _2919_ (.A1(_1380_),
    .A2(_1395_),
    .B1(_1396_),
    .Y(_0814_));
 sky130_fd_sc_hd__and3_1 _2920_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[40].S.IN1_L2 ),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1397_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2b_1 _2922_ (.A_N(_0816_),
    .B(_1396_),
    .Y(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_1398_),
    .X(_0815_));
 sky130_fd_sc_hd__a22oi_2 _2924_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[81].S.IN1_L5 ),
    .B1(_1375_),
    .B2(\stage_gen[1].mux_gen[81].S.IN1_L3 ),
    .Y(_1399_));
 sky130_fd_sc_hd__and3_1 _2925_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[40].S.IN1_L4 ),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _2926_ (.A(_1400_),
    .X(_0818_));
 sky130_fd_sc_hd__o21bai_1 _2927_ (.A1(_1366_),
    .A2(_1399_),
    .B1_N(_0818_),
    .Y(_0817_));
 sky130_fd_sc_hd__a22oi_1 _2928_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[82].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[82].S.IN1_L3 ),
    .Y(_1401_));
 sky130_fd_sc_hd__nand2_1 _2929_ (.A(_1388_),
    .B(\stage_gen[2].mux_gen[41].S.IN1_L1 ),
    .Y(_1402_));
 sky130_fd_sc_hd__o21ai_1 _2930_ (.A1(_1380_),
    .A2(_1401_),
    .B1(_1402_),
    .Y(_0819_));
 sky130_fd_sc_hd__and3_1 _2931_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[41].S.IN1_L2 ),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _2932_ (.A(_1403_),
    .X(_0821_));
 sky130_fd_sc_hd__nand2b_1 _2933_ (.A_N(_0821_),
    .B(_1402_),
    .Y(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _2934_ (.A(_1404_),
    .X(_0820_));
 sky130_fd_sc_hd__clkbuf_4 _2935_ (.A(_1369_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_4 _2936_ (.A(_1374_),
    .X(_1406_));
 sky130_fd_sc_hd__a22oi_1 _2937_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[83].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[83].S.IN1_L3 ),
    .Y(_1407_));
 sky130_fd_sc_hd__and3_1 _2938_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[41].S.IN1_L4 ),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1408_),
    .X(_0823_));
 sky130_fd_sc_hd__o21bai_1 _2940_ (.A1(_1366_),
    .A2(_1407_),
    .B1_N(_0823_),
    .Y(_0822_));
 sky130_fd_sc_hd__a22oi_1 _2941_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[84].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[84].S.IN1_L3 ),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2_1 _2942_ (.A(_1388_),
    .B(\stage_gen[2].mux_gen[42].S.IN1_L1 ),
    .Y(_1410_));
 sky130_fd_sc_hd__o21ai_1 _2943_ (.A1(_1380_),
    .A2(_1409_),
    .B1(_1410_),
    .Y(_0824_));
 sky130_fd_sc_hd__and3_1 _2944_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[42].S.IN1_L2 ),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_1411_),
    .X(_0826_));
 sky130_fd_sc_hd__nand2b_1 _2946_ (.A_N(_0826_),
    .B(_1410_),
    .Y(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _2947_ (.A(_1412_),
    .X(_0825_));
 sky130_fd_sc_hd__a22oi_2 _2948_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[85].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[85].S.IN1_L3 ),
    .Y(_1413_));
 sky130_fd_sc_hd__and3_1 _2949_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[42].S.IN1_L4 ),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1414_),
    .X(_0828_));
 sky130_fd_sc_hd__o21bai_1 _2951_ (.A1(_1366_),
    .A2(_1413_),
    .B1_N(_0828_),
    .Y(_0827_));
 sky130_fd_sc_hd__a22oi_1 _2952_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[86].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[86].S.IN1_L3 ),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_1 _2953_ (.A(_1388_),
    .B(\stage_gen[2].mux_gen[43].S.IN1_L1 ),
    .Y(_1416_));
 sky130_fd_sc_hd__o21ai_1 _2954_ (.A1(_1380_),
    .A2(_1415_),
    .B1(_1416_),
    .Y(_0829_));
 sky130_fd_sc_hd__and3_1 _2955_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[43].S.IN1_L2 ),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1417_),
    .X(_0831_));
 sky130_fd_sc_hd__nand2b_1 _2957_ (.A_N(_0831_),
    .B(_1416_),
    .Y(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1418_),
    .X(_0830_));
 sky130_fd_sc_hd__a22oi_1 _2959_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[87].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[87].S.IN1_L3 ),
    .Y(_1419_));
 sky130_fd_sc_hd__and3_1 _2960_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[43].S.IN1_L4 ),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1420_),
    .X(_0833_));
 sky130_fd_sc_hd__o21bai_1 _2962_ (.A1(_1366_),
    .A2(_1419_),
    .B1_N(_0833_),
    .Y(_0832_));
 sky130_fd_sc_hd__buf_4 _2963_ (.A(_1363_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_4 _2964_ (.A(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__a22oi_1 _2965_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[88].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[88].S.IN1_L3 ),
    .Y(_1423_));
 sky130_fd_sc_hd__buf_4 _2966_ (.A(_1387_),
    .X(_1424_));
 sky130_fd_sc_hd__nand2_1 _2967_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[44].S.IN1_L1 ),
    .Y(_1425_));
 sky130_fd_sc_hd__o21ai_1 _2968_ (.A1(_1422_),
    .A2(_1423_),
    .B1(_1425_),
    .Y(_0834_));
 sky130_fd_sc_hd__and3_1 _2969_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[44].S.IN1_L2 ),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1426_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2b_1 _2971_ (.A_N(_0836_),
    .B(_1425_),
    .Y(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1427_),
    .X(_0835_));
 sky130_fd_sc_hd__a22oi_2 _2973_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[89].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[89].S.IN1_L3 ),
    .Y(_1428_));
 sky130_fd_sc_hd__and3_1 _2974_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[44].S.IN1_L4 ),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _2975_ (.A(_1429_),
    .X(_0838_));
 sky130_fd_sc_hd__o21bai_1 _2976_ (.A1(_1366_),
    .A2(_1428_),
    .B1_N(_0838_),
    .Y(_0837_));
 sky130_fd_sc_hd__a22oi_1 _2977_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[90].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[90].S.IN1_L3 ),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _2978_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[45].S.IN1_L1 ),
    .Y(_1431_));
 sky130_fd_sc_hd__o21ai_1 _2979_ (.A1(_1422_),
    .A2(_1430_),
    .B1(_1431_),
    .Y(_0839_));
 sky130_fd_sc_hd__and3_1 _2980_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[45].S.IN1_L2 ),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1432_),
    .X(_0841_));
 sky130_fd_sc_hd__nand2b_1 _2982_ (.A_N(_0841_),
    .B(_1431_),
    .Y(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1433_),
    .X(_0840_));
 sky130_fd_sc_hd__a22oi_1 _2984_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[91].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[91].S.IN1_L3 ),
    .Y(_1434_));
 sky130_fd_sc_hd__and3_1 _2985_ (.A(_1364_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[45].S.IN1_L4 ),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_1435_),
    .X(_0843_));
 sky130_fd_sc_hd__o21bai_1 _2987_ (.A1(_1366_),
    .A2(_1434_),
    .B1_N(_0843_),
    .Y(_0842_));
 sky130_fd_sc_hd__a22oi_1 _2988_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[92].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[92].S.IN1_L3 ),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _2989_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[46].S.IN1_L1 ),
    .Y(_1437_));
 sky130_fd_sc_hd__o21ai_1 _2990_ (.A1(_1422_),
    .A2(_1436_),
    .B1(_1437_),
    .Y(_0844_));
 sky130_fd_sc_hd__and3_1 _2991_ (.A(_1359_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[46].S.IN1_L2 ),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _2992_ (.A(_1438_),
    .X(_0846_));
 sky130_fd_sc_hd__nand2b_1 _2993_ (.A_N(_0846_),
    .B(_1437_),
    .Y(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _2994_ (.A(_1439_),
    .X(_0845_));
 sky130_fd_sc_hd__a22oi_1 _2995_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[93].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[93].S.IN1_L3 ),
    .Y(_1440_));
 sky130_fd_sc_hd__buf_2 _2996_ (.A(_1363_),
    .X(_1441_));
 sky130_fd_sc_hd__and3_1 _2997_ (.A(_1441_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[46].S.IN1_L4 ),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_1442_),
    .X(_0848_));
 sky130_fd_sc_hd__o21bai_1 _2999_ (.A1(_1366_),
    .A2(_1440_),
    .B1_N(_0848_),
    .Y(_0847_));
 sky130_fd_sc_hd__a22oi_1 _3000_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[94].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[94].S.IN1_L3 ),
    .Y(_1443_));
 sky130_fd_sc_hd__nand2_1 _3001_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[47].S.IN1_L1 ),
    .Y(_1444_));
 sky130_fd_sc_hd__o21ai_1 _3002_ (.A1(_1422_),
    .A2(_1443_),
    .B1(_1444_),
    .Y(_0849_));
 sky130_fd_sc_hd__buf_4 _3003_ (.A(_1358_),
    .X(_1445_));
 sky130_fd_sc_hd__buf_2 _3004_ (.A(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__and3_1 _3005_ (.A(_1446_),
    .B(_1390_),
    .C(\stage_gen[2].mux_gen[47].S.IN1_L2 ),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1447_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2b_1 _3007_ (.A_N(_0851_),
    .B(_1444_),
    .Y(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _3008_ (.A(_1448_),
    .X(_0850_));
 sky130_fd_sc_hd__a22oi_1 _3009_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[95].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[95].S.IN1_L3 ),
    .Y(_1449_));
 sky130_fd_sc_hd__and3_1 _3010_ (.A(_1441_),
    .B(_1378_),
    .C(\stage_gen[2].mux_gen[47].S.IN1_L4 ),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_1450_),
    .X(_0853_));
 sky130_fd_sc_hd__o21bai_1 _3012_ (.A1(_1366_),
    .A2(_1449_),
    .B1_N(_0853_),
    .Y(_0852_));
 sky130_fd_sc_hd__clkbuf_4 _3013_ (.A(_1369_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_4 _3014_ (.A(_1374_),
    .X(_1452_));
 sky130_fd_sc_hd__a22oi_1 _3015_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[96].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[96].S.IN1_L3 ),
    .Y(_1453_));
 sky130_fd_sc_hd__nand2_1 _3016_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[48].S.IN1_L1 ),
    .Y(_1454_));
 sky130_fd_sc_hd__o21ai_1 _3017_ (.A1(_1422_),
    .A2(_1453_),
    .B1(_1454_),
    .Y(_0854_));
 sky130_fd_sc_hd__clkbuf_4 _3018_ (.A(_1360_),
    .X(_1455_));
 sky130_fd_sc_hd__and3_1 _3019_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[48].S.IN1_L2 ),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _3020_ (.A(_1456_),
    .X(_0856_));
 sky130_fd_sc_hd__nand2b_1 _3021_ (.A_N(_0856_),
    .B(_1454_),
    .Y(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3022_ (.A(_1457_),
    .X(_0855_));
 sky130_fd_sc_hd__buf_2 _3023_ (.A(_1421_),
    .X(_1458_));
 sky130_fd_sc_hd__a22oi_1 _3024_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[97].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[97].S.IN1_L3 ),
    .Y(_1459_));
 sky130_fd_sc_hd__clkbuf_2 _3025_ (.A(_1377_),
    .X(_1460_));
 sky130_fd_sc_hd__and3_1 _3026_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[48].S.IN1_L4 ),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_1461_),
    .X(_0858_));
 sky130_fd_sc_hd__o21bai_1 _3028_ (.A1(_1458_),
    .A2(_1459_),
    .B1_N(_0858_),
    .Y(_0857_));
 sky130_fd_sc_hd__a22oi_1 _3029_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[98].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[98].S.IN1_L3 ),
    .Y(_1462_));
 sky130_fd_sc_hd__nand2_1 _3030_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[49].S.IN1_L1 ),
    .Y(_1463_));
 sky130_fd_sc_hd__o21ai_1 _3031_ (.A1(_1422_),
    .A2(_1462_),
    .B1(_1463_),
    .Y(_0859_));
 sky130_fd_sc_hd__and3_1 _3032_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[49].S.IN1_L2 ),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1464_),
    .X(_0861_));
 sky130_fd_sc_hd__nand2b_1 _3034_ (.A_N(_0861_),
    .B(_1463_),
    .Y(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1465_),
    .X(_0860_));
 sky130_fd_sc_hd__a22oi_1 _3036_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[99].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[99].S.IN1_L3 ),
    .Y(_1466_));
 sky130_fd_sc_hd__and3_1 _3037_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[49].S.IN1_L4 ),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3038_ (.A(_1467_),
    .X(_0863_));
 sky130_fd_sc_hd__o21bai_1 _3039_ (.A1(_1458_),
    .A2(_1466_),
    .B1_N(_0863_),
    .Y(_0862_));
 sky130_fd_sc_hd__a22oi_1 _3040_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[100].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[100].S.IN1_L3 ),
    .Y(_1468_));
 sky130_fd_sc_hd__nand2_1 _3041_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[50].S.IN1_L1 ),
    .Y(_1469_));
 sky130_fd_sc_hd__o21ai_1 _3042_ (.A1(_1422_),
    .A2(_1468_),
    .B1(_1469_),
    .Y(_0869_));
 sky130_fd_sc_hd__and3_1 _3043_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[50].S.IN1_L2 ),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1470_),
    .X(_0871_));
 sky130_fd_sc_hd__nand2b_1 _3045_ (.A_N(_0871_),
    .B(_1469_),
    .Y(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1471_),
    .X(_0870_));
 sky130_fd_sc_hd__a22oi_1 _3047_ (.A1(_1405_),
    .A2(\stage_gen[1].mux_gen[101].S.IN1_L5 ),
    .B1(_1406_),
    .B2(\stage_gen[1].mux_gen[101].S.IN1_L3 ),
    .Y(_1472_));
 sky130_fd_sc_hd__and3_1 _3048_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[50].S.IN1_L4 ),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3049_ (.A(_1473_),
    .X(_0873_));
 sky130_fd_sc_hd__o21bai_1 _3050_ (.A1(_1458_),
    .A2(_1472_),
    .B1_N(_0873_),
    .Y(_0872_));
 sky130_fd_sc_hd__a22oi_1 _3051_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[102].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[102].S.IN1_L3 ),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _3052_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[51].S.IN1_L1 ),
    .Y(_1475_));
 sky130_fd_sc_hd__o21ai_1 _3053_ (.A1(_1422_),
    .A2(_1474_),
    .B1(_1475_),
    .Y(_0874_));
 sky130_fd_sc_hd__and3_1 _3054_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[51].S.IN1_L2 ),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1476_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2b_1 _3056_ (.A_N(_0876_),
    .B(_1475_),
    .Y(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3057_ (.A(_1477_),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _3058_ (.A(_1369_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_4 _3059_ (.A(_1374_),
    .X(_1479_));
 sky130_fd_sc_hd__a22oi_1 _3060_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[103].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[103].S.IN1_L3 ),
    .Y(_1480_));
 sky130_fd_sc_hd__and3_1 _3061_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[51].S.IN1_L4 ),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1481_),
    .X(_0878_));
 sky130_fd_sc_hd__o21bai_1 _3063_ (.A1(_1458_),
    .A2(_1480_),
    .B1_N(_0878_),
    .Y(_0877_));
 sky130_fd_sc_hd__a22oi_1 _3064_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[104].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[104].S.IN1_L3 ),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _3065_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[52].S.IN1_L1 ),
    .Y(_1483_));
 sky130_fd_sc_hd__o21ai_1 _3066_ (.A1(_1422_),
    .A2(_1482_),
    .B1(_1483_),
    .Y(_0879_));
 sky130_fd_sc_hd__and3_1 _3067_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[52].S.IN1_L2 ),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3068_ (.A(_1484_),
    .X(_0881_));
 sky130_fd_sc_hd__nand2b_1 _3069_ (.A_N(_0881_),
    .B(_1483_),
    .Y(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3070_ (.A(_1485_),
    .X(_0880_));
 sky130_fd_sc_hd__a22oi_1 _3071_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[105].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[105].S.IN1_L3 ),
    .Y(_1486_));
 sky130_fd_sc_hd__and3_1 _3072_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[52].S.IN1_L4 ),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1487_),
    .X(_0883_));
 sky130_fd_sc_hd__o21bai_1 _3074_ (.A1(_1458_),
    .A2(_1486_),
    .B1_N(_0883_),
    .Y(_0882_));
 sky130_fd_sc_hd__a22oi_1 _3075_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[106].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[106].S.IN1_L3 ),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(_1424_),
    .B(\stage_gen[2].mux_gen[53].S.IN1_L1 ),
    .Y(_1489_));
 sky130_fd_sc_hd__o21ai_1 _3077_ (.A1(_1422_),
    .A2(_1488_),
    .B1(_1489_),
    .Y(_0884_));
 sky130_fd_sc_hd__and3_1 _3078_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[53].S.IN1_L2 ),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3079_ (.A(_1490_),
    .X(_0886_));
 sky130_fd_sc_hd__nand2b_1 _3080_ (.A_N(_0886_),
    .B(_1489_),
    .Y(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3081_ (.A(_1491_),
    .X(_0885_));
 sky130_fd_sc_hd__a22oi_1 _3082_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[107].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[107].S.IN1_L3 ),
    .Y(_1492_));
 sky130_fd_sc_hd__and3_1 _3083_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[53].S.IN1_L4 ),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1493_),
    .X(_0888_));
 sky130_fd_sc_hd__o21bai_1 _3085_ (.A1(_1458_),
    .A2(_1492_),
    .B1_N(_0888_),
    .Y(_0887_));
 sky130_fd_sc_hd__clkbuf_4 _3086_ (.A(_1421_),
    .X(_1494_));
 sky130_fd_sc_hd__a22oi_1 _3087_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[108].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[108].S.IN1_L3 ),
    .Y(_1495_));
 sky130_fd_sc_hd__clkbuf_4 _3088_ (.A(_1387_),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _3089_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[54].S.IN1_L1 ),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_1 _3090_ (.A1(_1494_),
    .A2(_1495_),
    .B1(_1497_),
    .Y(_0889_));
 sky130_fd_sc_hd__and3_1 _3091_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[54].S.IN1_L2 ),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3092_ (.A(_1498_),
    .X(_0891_));
 sky130_fd_sc_hd__nand2b_1 _3093_ (.A_N(_0891_),
    .B(_1497_),
    .Y(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1499_),
    .X(_0890_));
 sky130_fd_sc_hd__a22oi_1 _3095_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[109].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[109].S.IN1_L3 ),
    .Y(_1500_));
 sky130_fd_sc_hd__and3_1 _3096_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[54].S.IN1_L4 ),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3097_ (.A(_1501_),
    .X(_0893_));
 sky130_fd_sc_hd__o21bai_1 _3098_ (.A1(_1458_),
    .A2(_1500_),
    .B1_N(_0893_),
    .Y(_0892_));
 sky130_fd_sc_hd__a22oi_1 _3099_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[110].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[110].S.IN1_L3 ),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _3100_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[55].S.IN1_L1 ),
    .Y(_1503_));
 sky130_fd_sc_hd__o21ai_1 _3101_ (.A1(_1494_),
    .A2(_1502_),
    .B1(_1503_),
    .Y(_0894_));
 sky130_fd_sc_hd__and3_1 _3102_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[55].S.IN1_L2 ),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3103_ (.A(_1504_),
    .X(_0896_));
 sky130_fd_sc_hd__nand2b_1 _3104_ (.A_N(_0896_),
    .B(_1503_),
    .Y(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3105_ (.A(_1505_),
    .X(_0895_));
 sky130_fd_sc_hd__a22oi_2 _3106_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[111].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[111].S.IN1_L3 ),
    .Y(_1506_));
 sky130_fd_sc_hd__and3_1 _3107_ (.A(_1441_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[55].S.IN1_L4 ),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1507_),
    .X(_0898_));
 sky130_fd_sc_hd__o21bai_1 _3109_ (.A1(_1458_),
    .A2(_1506_),
    .B1_N(_0898_),
    .Y(_0897_));
 sky130_fd_sc_hd__a22oi_1 _3110_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[112].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[112].S.IN1_L3 ),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2_1 _3111_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[56].S.IN1_L1 ),
    .Y(_1509_));
 sky130_fd_sc_hd__o21ai_1 _3112_ (.A1(_1494_),
    .A2(_1508_),
    .B1(_1509_),
    .Y(_0899_));
 sky130_fd_sc_hd__and3_1 _3113_ (.A(_1446_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[56].S.IN1_L2 ),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3114_ (.A(_1510_),
    .X(_0901_));
 sky130_fd_sc_hd__nand2b_1 _3115_ (.A_N(_0901_),
    .B(_1509_),
    .Y(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3116_ (.A(_1511_),
    .X(_0900_));
 sky130_fd_sc_hd__a22oi_1 _3117_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[113].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[113].S.IN1_L3 ),
    .Y(_1512_));
 sky130_fd_sc_hd__buf_2 _3118_ (.A(_1363_),
    .X(_1513_));
 sky130_fd_sc_hd__and3_1 _3119_ (.A(_1513_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[56].S.IN1_L4 ),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1514_),
    .X(_0903_));
 sky130_fd_sc_hd__o21bai_1 _3121_ (.A1(_1458_),
    .A2(_1512_),
    .B1_N(_0903_),
    .Y(_0902_));
 sky130_fd_sc_hd__a22oi_1 _3122_ (.A1(_1451_),
    .A2(\stage_gen[1].mux_gen[114].S.IN1_L5 ),
    .B1(_1452_),
    .B2(\stage_gen[1].mux_gen[114].S.IN1_L3 ),
    .Y(_1515_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[57].S.IN1_L1 ),
    .Y(_1516_));
 sky130_fd_sc_hd__o21ai_1 _3124_ (.A1(_1494_),
    .A2(_1515_),
    .B1(_1516_),
    .Y(_0904_));
 sky130_fd_sc_hd__buf_2 _3125_ (.A(_1445_),
    .X(_1517_));
 sky130_fd_sc_hd__and3_1 _3126_ (.A(_1517_),
    .B(_1455_),
    .C(\stage_gen[2].mux_gen[57].S.IN1_L2 ),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3127_ (.A(_1518_),
    .X(_0906_));
 sky130_fd_sc_hd__nand2b_1 _3128_ (.A_N(_0906_),
    .B(_1516_),
    .Y(_1519_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_1519_),
    .X(_0905_));
 sky130_fd_sc_hd__a22oi_2 _3130_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[115].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[115].S.IN1_L3 ),
    .Y(_1520_));
 sky130_fd_sc_hd__and3_1 _3131_ (.A(_1513_),
    .B(_1460_),
    .C(\stage_gen[2].mux_gen[57].S.IN1_L4 ),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3132_ (.A(_1521_),
    .X(_0908_));
 sky130_fd_sc_hd__o21bai_1 _3133_ (.A1(_1458_),
    .A2(_1520_),
    .B1_N(_0908_),
    .Y(_0907_));
 sky130_fd_sc_hd__clkbuf_4 _3134_ (.A(_1369_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_4 _3135_ (.A(_1374_),
    .X(_1523_));
 sky130_fd_sc_hd__a22oi_1 _3136_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[116].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[116].S.IN1_L3 ),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_1 _3137_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[58].S.IN1_L1 ),
    .Y(_1525_));
 sky130_fd_sc_hd__o21ai_1 _3138_ (.A1(_1494_),
    .A2(_1524_),
    .B1(_1525_),
    .Y(_0909_));
 sky130_fd_sc_hd__clkbuf_4 _3139_ (.A(_1360_),
    .X(_1526_));
 sky130_fd_sc_hd__and3_1 _3140_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[58].S.IN1_L2 ),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3141_ (.A(_1527_),
    .X(_0911_));
 sky130_fd_sc_hd__nand2b_1 _3142_ (.A_N(_0911_),
    .B(_1525_),
    .Y(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1528_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_4 _3144_ (.A(_1421_),
    .X(_1529_));
 sky130_fd_sc_hd__a22oi_1 _3145_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[117].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[117].S.IN1_L3 ),
    .Y(_1530_));
 sky130_fd_sc_hd__buf_2 _3146_ (.A(_1377_),
    .X(_1531_));
 sky130_fd_sc_hd__and3_1 _3147_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[58].S.IN1_L4 ),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3148_ (.A(_1532_),
    .X(_0913_));
 sky130_fd_sc_hd__o21bai_1 _3149_ (.A1(_1529_),
    .A2(_1530_),
    .B1_N(_0913_),
    .Y(_0912_));
 sky130_fd_sc_hd__a22oi_1 _3150_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[118].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[118].S.IN1_L3 ),
    .Y(_1533_));
 sky130_fd_sc_hd__nand2_1 _3151_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[59].S.IN1_L1 ),
    .Y(_1534_));
 sky130_fd_sc_hd__o21ai_1 _3152_ (.A1(_1494_),
    .A2(_1533_),
    .B1(_1534_),
    .Y(_0914_));
 sky130_fd_sc_hd__and3_1 _3153_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[59].S.IN1_L2 ),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1535_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2b_1 _3155_ (.A_N(_0916_),
    .B(_1534_),
    .Y(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1536_),
    .X(_0915_));
 sky130_fd_sc_hd__a22oi_1 _3157_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[119].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[119].S.IN1_L3 ),
    .Y(_1537_));
 sky130_fd_sc_hd__and3_1 _3158_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[59].S.IN1_L4 ),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1538_),
    .X(_0918_));
 sky130_fd_sc_hd__o21bai_1 _3160_ (.A1(_1529_),
    .A2(_1537_),
    .B1_N(_0918_),
    .Y(_0917_));
 sky130_fd_sc_hd__a22oi_1 _3161_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[120].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[120].S.IN1_L3 ),
    .Y(_1539_));
 sky130_fd_sc_hd__nand2_1 _3162_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[60].S.IN1_L1 ),
    .Y(_1540_));
 sky130_fd_sc_hd__o21ai_1 _3163_ (.A1(_1494_),
    .A2(_1539_),
    .B1(_1540_),
    .Y(_0924_));
 sky130_fd_sc_hd__and3_1 _3164_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[60].S.IN1_L2 ),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3165_ (.A(_1541_),
    .X(_0926_));
 sky130_fd_sc_hd__nand2b_1 _3166_ (.A_N(_0926_),
    .B(_1540_),
    .Y(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3167_ (.A(_1542_),
    .X(_0925_));
 sky130_fd_sc_hd__a22oi_1 _3168_ (.A1(_1478_),
    .A2(\stage_gen[1].mux_gen[121].S.IN1_L5 ),
    .B1(_1479_),
    .B2(\stage_gen[1].mux_gen[121].S.IN1_L3 ),
    .Y(_1543_));
 sky130_fd_sc_hd__and3_1 _3169_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[60].S.IN1_L4 ),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1544_),
    .X(_0928_));
 sky130_fd_sc_hd__o21bai_1 _3171_ (.A1(_1529_),
    .A2(_1543_),
    .B1_N(_0928_),
    .Y(_0927_));
 sky130_fd_sc_hd__a22oi_1 _3172_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[122].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[122].S.IN1_L3 ),
    .Y(_1545_));
 sky130_fd_sc_hd__nand2_1 _3173_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[61].S.IN1_L1 ),
    .Y(_1546_));
 sky130_fd_sc_hd__o21ai_1 _3174_ (.A1(_1494_),
    .A2(_1545_),
    .B1(_1546_),
    .Y(_0929_));
 sky130_fd_sc_hd__and3_1 _3175_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[61].S.IN1_L2 ),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1547_),
    .X(_0931_));
 sky130_fd_sc_hd__nand2b_1 _3177_ (.A_N(_0931_),
    .B(_1546_),
    .Y(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1548_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_4 _3179_ (.A(_1369_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_4 _3180_ (.A(_1374_),
    .X(_1550_));
 sky130_fd_sc_hd__a22oi_1 _3181_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[123].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[123].S.IN1_L3 ),
    .Y(_1551_));
 sky130_fd_sc_hd__and3_1 _3182_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[61].S.IN1_L4 ),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1552_),
    .X(_0933_));
 sky130_fd_sc_hd__o21bai_1 _3184_ (.A1(_1529_),
    .A2(_1551_),
    .B1_N(_0933_),
    .Y(_0932_));
 sky130_fd_sc_hd__a22oi_1 _3185_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[124].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[124].S.IN1_L3 ),
    .Y(_1553_));
 sky130_fd_sc_hd__nand2_1 _3186_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[62].S.IN1_L1 ),
    .Y(_1554_));
 sky130_fd_sc_hd__o21ai_1 _3187_ (.A1(_1494_),
    .A2(_1553_),
    .B1(_1554_),
    .Y(_0934_));
 sky130_fd_sc_hd__and3_1 _3188_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[62].S.IN1_L2 ),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1555_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2b_1 _3190_ (.A_N(_0936_),
    .B(_1554_),
    .Y(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1556_),
    .X(_0935_));
 sky130_fd_sc_hd__a22oi_1 _3192_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[125].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[125].S.IN1_L3 ),
    .Y(_1557_));
 sky130_fd_sc_hd__and3_1 _3193_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[62].S.IN1_L4 ),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1558_),
    .X(_0938_));
 sky130_fd_sc_hd__o21bai_1 _3195_ (.A1(_1529_),
    .A2(_1557_),
    .B1_N(_0938_),
    .Y(_0937_));
 sky130_fd_sc_hd__a22oi_1 _3196_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[126].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[126].S.IN1_L3 ),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _3197_ (.A(_1496_),
    .B(\stage_gen[2].mux_gen[63].S.IN1_L1 ),
    .Y(_1560_));
 sky130_fd_sc_hd__o21ai_1 _3198_ (.A1(_1494_),
    .A2(_1559_),
    .B1(_1560_),
    .Y(_0939_));
 sky130_fd_sc_hd__and3_1 _3199_ (.A(_1517_),
    .B(_1526_),
    .C(\stage_gen[2].mux_gen[63].S.IN1_L2 ),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3200_ (.A(_1561_),
    .X(_0941_));
 sky130_fd_sc_hd__nand2b_1 _3201_ (.A_N(_0941_),
    .B(_1560_),
    .Y(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3202_ (.A(_1562_),
    .X(_0940_));
 sky130_fd_sc_hd__a22oi_1 _3203_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[127].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[127].S.IN1_L3 ),
    .Y(_1563_));
 sky130_fd_sc_hd__and3_1 _3204_ (.A(_1513_),
    .B(_1531_),
    .C(\stage_gen[2].mux_gen[63].S.IN1_L4 ),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1564_),
    .X(_0943_));
 sky130_fd_sc_hd__o21bai_1 _3206_ (.A1(_1529_),
    .A2(_1563_),
    .B1_N(_0943_),
    .Y(_0942_));
 sky130_fd_sc_hd__clkbuf_2 _3207_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .X(_1565_));
 sky130_fd_sc_hd__buf_4 _3208_ (.A(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__buf_6 _3209_ (.A(_1387_),
    .X(_1567_));
 sky130_fd_sc_hd__nand2_1 _3210_ (.A(_1358_),
    .B(_1384_),
    .Y(_1568_));
 sky130_fd_sc_hd__inv_2 _3211_ (.A(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__buf_4 _3212_ (.A(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__buf_6 _3213_ (.A(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__a22oi_2 _3214_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[0].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[0].S.IN1_L3 ),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _3215_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .B(net257),
    .Y(_1573_));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__clkbuf_4 _3217_ (.A(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__buf_4 _3218_ (.A(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nand2_1 _3219_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[0].S.IN1_L1 ),
    .Y(_1577_));
 sky130_fd_sc_hd__o21ai_1 _3220_ (.A1(_1566_),
    .A2(_1572_),
    .B1(_1577_),
    .Y(_0964_));
 sky130_fd_sc_hd__inv_2 _3221_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .Y(_1578_));
 sky130_fd_sc_hd__buf_2 _3222_ (.A(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__and3_1 _3223_ (.A(_1579_),
    .B(_1526_),
    .C(\stage_gen[3].mux_gen[0].S.IN1_L2 ),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1580_),
    .X(_0966_));
 sky130_fd_sc_hd__nand2b_1 _3225_ (.A_N(_0966_),
    .B(_1577_),
    .Y(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1581_),
    .X(_0965_));
 sky130_fd_sc_hd__buf_4 _3227_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_4 _3228_ (.A(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_2 _3229_ (.A(_1387_),
    .X(_0647_));
 sky130_fd_sc_hd__buf_6 _3230_ (.A(_1570_),
    .X(_0648_));
 sky130_fd_sc_hd__a22oi_2 _3231_ (.A1(net414),
    .A2(\stage_gen[2].mux_gen[1].S.IN1_L5 ),
    .B1(net311),
    .B2(\stage_gen[2].mux_gen[1].S.IN1_L3 ),
    .Y(_1584_));
 sky130_fd_sc_hd__and3_1 _3232_ (.A(_1565_),
    .B(_1531_),
    .C(\stage_gen[3].mux_gen[0].S.IN1_L4 ),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3233_ (.A(_1585_),
    .X(_0968_));
 sky130_fd_sc_hd__o21bai_1 _3234_ (.A1(_1583_),
    .A2(_1584_),
    .B1_N(_0968_),
    .Y(_0967_));
 sky130_fd_sc_hd__a22oi_2 _3235_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[2].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[2].S.IN1_L3 ),
    .Y(_1586_));
 sky130_fd_sc_hd__nand2_1 _3236_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[1].S.IN1_L1 ),
    .Y(_1587_));
 sky130_fd_sc_hd__o21ai_1 _3237_ (.A1(_1566_),
    .A2(_1586_),
    .B1(_1587_),
    .Y(_1021_));
 sky130_fd_sc_hd__and3_1 _3238_ (.A(_1579_),
    .B(_1526_),
    .C(\stage_gen[3].mux_gen[1].S.IN1_L2 ),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3239_ (.A(_1588_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2b_1 _3240_ (.A_N(_1023_),
    .B(_1587_),
    .Y(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_1589_),
    .X(_1022_));
 sky130_fd_sc_hd__a22oi_2 _3242_ (.A1(net415),
    .A2(\stage_gen[2].mux_gen[3].S.IN1_L5 ),
    .B1(net310),
    .B2(\stage_gen[2].mux_gen[3].S.IN1_L3 ),
    .Y(_1590_));
 sky130_fd_sc_hd__and3_1 _3243_ (.A(_1565_),
    .B(_1531_),
    .C(\stage_gen[3].mux_gen[1].S.IN1_L4 ),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_1591_),
    .X(_1025_));
 sky130_fd_sc_hd__o21bai_1 _3245_ (.A1(_1583_),
    .A2(_1590_),
    .B1_N(_1025_),
    .Y(_1024_));
 sky130_fd_sc_hd__a22oi_4 _3246_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[4].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[4].S.IN1_L3 ),
    .Y(_1592_));
 sky130_fd_sc_hd__nand2_1 _3247_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[2].S.IN1_L1 ),
    .Y(_1593_));
 sky130_fd_sc_hd__o21ai_1 _3248_ (.A1(_1566_),
    .A2(_1592_),
    .B1(_1593_),
    .Y(_1076_));
 sky130_fd_sc_hd__and3_1 _3249_ (.A(_1579_),
    .B(_1526_),
    .C(\stage_gen[3].mux_gen[2].S.IN1_L2 ),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1594_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2b_1 _3251_ (.A_N(_1078_),
    .B(_1593_),
    .Y(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3252_ (.A(_1595_),
    .X(_1077_));
 sky130_fd_sc_hd__a22oi_2 _3253_ (.A1(net415),
    .A2(\stage_gen[2].mux_gen[5].S.IN1_L5 ),
    .B1(net310),
    .B2(\stage_gen[2].mux_gen[5].S.IN1_L3 ),
    .Y(_1596_));
 sky130_fd_sc_hd__and3_1 _3254_ (.A(_1565_),
    .B(_1531_),
    .C(\stage_gen[3].mux_gen[2].S.IN1_L4 ),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1597_),
    .X(_1080_));
 sky130_fd_sc_hd__o21bai_1 _3256_ (.A1(_1583_),
    .A2(_1596_),
    .B1_N(_1080_),
    .Y(_1079_));
 sky130_fd_sc_hd__a22oi_2 _3257_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[6].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[6].S.IN1_L3 ),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _3258_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[3].S.IN1_L1 ),
    .Y(_1599_));
 sky130_fd_sc_hd__o21ai_1 _3259_ (.A1(_1566_),
    .A2(_1598_),
    .B1(_1599_),
    .Y(_1091_));
 sky130_fd_sc_hd__and3_1 _3260_ (.A(_1579_),
    .B(_1526_),
    .C(\stage_gen[3].mux_gen[3].S.IN1_L2 ),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1600_),
    .X(_1093_));
 sky130_fd_sc_hd__nand2b_1 _3262_ (.A_N(_1093_),
    .B(_1599_),
    .Y(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3263_ (.A(_1601_),
    .X(_1092_));
 sky130_fd_sc_hd__a22oi_4 _3264_ (.A1(net410),
    .A2(\stage_gen[2].mux_gen[7].S.IN1_L5 ),
    .B1(net308),
    .B2(\stage_gen[2].mux_gen[7].S.IN1_L3 ),
    .Y(_1602_));
 sky130_fd_sc_hd__and3_1 _3265_ (.A(_1565_),
    .B(_1531_),
    .C(\stage_gen[3].mux_gen[3].S.IN1_L4 ),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3266_ (.A(_1603_),
    .X(_1095_));
 sky130_fd_sc_hd__o21bai_1 _3267_ (.A1(_1583_),
    .A2(_1602_),
    .B1_N(_1095_),
    .Y(_1094_));
 sky130_fd_sc_hd__a22oi_4 _3268_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[8].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[8].S.IN1_L3 ),
    .Y(_1604_));
 sky130_fd_sc_hd__nand2_1 _3269_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[4].S.IN1_L1 ),
    .Y(_1605_));
 sky130_fd_sc_hd__o21ai_1 _3270_ (.A1(_1566_),
    .A2(_1604_),
    .B1(_1605_),
    .Y(_1096_));
 sky130_fd_sc_hd__clkbuf_4 _3271_ (.A(_1360_),
    .X(_1606_));
 sky130_fd_sc_hd__and3_1 _3272_ (.A(_1579_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[4].S.IN1_L2 ),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1607_),
    .X(_1098_));
 sky130_fd_sc_hd__nand2b_1 _3274_ (.A_N(_1098_),
    .B(_1605_),
    .Y(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3275_ (.A(_1608_),
    .X(_1097_));
 sky130_fd_sc_hd__a22oi_4 _3276_ (.A1(net412),
    .A2(\stage_gen[2].mux_gen[9].S.IN1_L5 ),
    .B1(net309),
    .B2(\stage_gen[2].mux_gen[9].S.IN1_L3 ),
    .Y(_1609_));
 sky130_fd_sc_hd__buf_2 _3277_ (.A(_1377_),
    .X(_1610_));
 sky130_fd_sc_hd__and3_1 _3278_ (.A(_1565_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[4].S.IN1_L4 ),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1611_),
    .X(_1100_));
 sky130_fd_sc_hd__o21bai_1 _3280_ (.A1(_1583_),
    .A2(_1609_),
    .B1_N(_1100_),
    .Y(_1099_));
 sky130_fd_sc_hd__a22oi_4 _3281_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[10].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[10].S.IN1_L3 ),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[5].S.IN1_L1 ),
    .Y(_1613_));
 sky130_fd_sc_hd__o21ai_1 _3283_ (.A1(_1566_),
    .A2(_1612_),
    .B1(_1613_),
    .Y(_1101_));
 sky130_fd_sc_hd__and3_1 _3284_ (.A(_1579_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[5].S.IN1_L2 ),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3285_ (.A(_1614_),
    .X(_1103_));
 sky130_fd_sc_hd__nand2b_1 _3286_ (.A_N(_1103_),
    .B(_1613_),
    .Y(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3287_ (.A(_1615_),
    .X(_1102_));
 sky130_fd_sc_hd__a22oi_4 _3288_ (.A1(net406),
    .A2(\stage_gen[2].mux_gen[11].S.IN1_L5 ),
    .B1(net305),
    .B2(\stage_gen[2].mux_gen[11].S.IN1_L3 ),
    .Y(_1616_));
 sky130_fd_sc_hd__and3_1 _3289_ (.A(_1565_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[5].S.IN1_L4 ),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3290_ (.A(_1617_),
    .X(_1105_));
 sky130_fd_sc_hd__o21bai_1 _3291_ (.A1(_1583_),
    .A2(_1616_),
    .B1_N(_1105_),
    .Y(_1104_));
 sky130_fd_sc_hd__a22oi_2 _3292_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[12].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[12].S.IN1_L3 ),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _3293_ (.A(_1576_),
    .B(\stage_gen[3].mux_gen[6].S.IN1_L1 ),
    .Y(_1619_));
 sky130_fd_sc_hd__o21ai_1 _3294_ (.A1(_1566_),
    .A2(_1618_),
    .B1(_1619_),
    .Y(_1106_));
 sky130_fd_sc_hd__and3_1 _3295_ (.A(_1579_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[6].S.IN1_L2 ),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3296_ (.A(_1620_),
    .X(_1108_));
 sky130_fd_sc_hd__nand2b_1 _3297_ (.A_N(_1108_),
    .B(_1619_),
    .Y(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3298_ (.A(_1621_),
    .X(_1107_));
 sky130_fd_sc_hd__a22oi_4 _3299_ (.A1(net405),
    .A2(\stage_gen[2].mux_gen[13].S.IN1_L5 ),
    .B1(net304),
    .B2(\stage_gen[2].mux_gen[13].S.IN1_L3 ),
    .Y(_1622_));
 sky130_fd_sc_hd__and3_1 _3300_ (.A(_1565_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[6].S.IN1_L4 ),
    .X(_1623_));
 sky130_fd_sc_hd__buf_6 _3301_ (.A(_1623_),
    .X(_1110_));
 sky130_fd_sc_hd__o21bai_1 _3302_ (.A1(_1583_),
    .A2(_1622_),
    .B1_N(_1110_),
    .Y(_1109_));
 sky130_fd_sc_hd__buf_2 _3303_ (.A(_1582_),
    .X(_1624_));
 sky130_fd_sc_hd__buf_6 _3304_ (.A(_1387_),
    .X(_1625_));
 sky130_fd_sc_hd__buf_6 _3305_ (.A(_1570_),
    .X(_1626_));
 sky130_fd_sc_hd__a22oi_4 _3306_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[14].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[14].S.IN1_L3 ),
    .Y(_1627_));
 sky130_fd_sc_hd__buf_2 _3307_ (.A(_1575_),
    .X(_1628_));
 sky130_fd_sc_hd__nand2_1 _3308_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[7].S.IN1_L1 ),
    .Y(_1629_));
 sky130_fd_sc_hd__o21ai_1 _3309_ (.A1(_1624_),
    .A2(_1627_),
    .B1(_1629_),
    .Y(_1111_));
 sky130_fd_sc_hd__and3_1 _3310_ (.A(_1579_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[7].S.IN1_L2 ),
    .X(_1630_));
 sky130_fd_sc_hd__clkbuf_1 _3311_ (.A(_1630_),
    .X(_1113_));
 sky130_fd_sc_hd__nand2b_1 _3312_ (.A_N(_1113_),
    .B(_1629_),
    .Y(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3313_ (.A(_1631_),
    .X(_1112_));
 sky130_fd_sc_hd__a22oi_4 _3314_ (.A1(net404),
    .A2(\stage_gen[2].mux_gen[15].S.IN1_L5 ),
    .B1(net304),
    .B2(\stage_gen[2].mux_gen[15].S.IN1_L3 ),
    .Y(_1632_));
 sky130_fd_sc_hd__and3_1 _3315_ (.A(_1565_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[7].S.IN1_L4 ),
    .X(_1633_));
 sky130_fd_sc_hd__buf_6 _3316_ (.A(_1633_),
    .X(_1115_));
 sky130_fd_sc_hd__o21bai_1 _3317_ (.A1(_1583_),
    .A2(_1632_),
    .B1_N(_1115_),
    .Y(_1114_));
 sky130_fd_sc_hd__a22oi_4 _3318_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[16].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[16].S.IN1_L3 ),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2_1 _3319_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[8].S.IN1_L1 ),
    .Y(_1635_));
 sky130_fd_sc_hd__o21ai_1 _3320_ (.A1(_1624_),
    .A2(_1634_),
    .B1(_1635_),
    .Y(_1116_));
 sky130_fd_sc_hd__buf_2 _3321_ (.A(_1578_),
    .X(_1636_));
 sky130_fd_sc_hd__and3_1 _3322_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[8].S.IN1_L2 ),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _3323_ (.A(_1637_),
    .X(_1118_));
 sky130_fd_sc_hd__nand2b_1 _3324_ (.A_N(_1118_),
    .B(_1635_),
    .Y(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1638_),
    .X(_1117_));
 sky130_fd_sc_hd__a22oi_4 _3326_ (.A1(net407),
    .A2(\stage_gen[2].mux_gen[17].S.IN1_L5 ),
    .B1(net306),
    .B2(\stage_gen[2].mux_gen[17].S.IN1_L3 ),
    .Y(_1639_));
 sky130_fd_sc_hd__and3_1 _3327_ (.A(_1565_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[8].S.IN1_L4 ),
    .X(_1640_));
 sky130_fd_sc_hd__buf_6 _3328_ (.A(_1640_),
    .X(_1120_));
 sky130_fd_sc_hd__o21bai_1 _3329_ (.A1(_1583_),
    .A2(_1639_),
    .B1_N(_1120_),
    .Y(_1119_));
 sky130_fd_sc_hd__a22oi_4 _3330_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[18].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[18].S.IN1_L3 ),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[9].S.IN1_L1 ),
    .Y(_1642_));
 sky130_fd_sc_hd__o21ai_1 _3332_ (.A1(_1624_),
    .A2(_1641_),
    .B1(_1642_),
    .Y(_1121_));
 sky130_fd_sc_hd__and3_1 _3333_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[9].S.IN1_L2 ),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _3334_ (.A(_1643_),
    .X(_1123_));
 sky130_fd_sc_hd__nand2b_1 _3335_ (.A_N(_1123_),
    .B(_1642_),
    .Y(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3336_ (.A(_1644_),
    .X(_1122_));
 sky130_fd_sc_hd__buf_4 _3337_ (.A(_1386_),
    .X(_1645_));
 sky130_fd_sc_hd__buf_6 _3338_ (.A(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__buf_6 _3339_ (.A(_1570_),
    .X(_1647_));
 sky130_fd_sc_hd__a22oi_4 _3340_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[19].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[19].S.IN1_L3 ),
    .Y(_1648_));
 sky130_fd_sc_hd__clkbuf_2 _3341_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .X(_1649_));
 sky130_fd_sc_hd__and3_1 _3342_ (.A(_1649_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[9].S.IN1_L4 ),
    .X(_1650_));
 sky130_fd_sc_hd__buf_6 _3343_ (.A(_1650_),
    .X(_1125_));
 sky130_fd_sc_hd__o21bai_1 _3344_ (.A1(_1583_),
    .A2(_1648_),
    .B1_N(_1125_),
    .Y(_1124_));
 sky130_fd_sc_hd__a22oi_4 _3345_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[20].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[20].S.IN1_L3 ),
    .Y(_1651_));
 sky130_fd_sc_hd__nand2_1 _3346_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[10].S.IN1_L1 ),
    .Y(_1652_));
 sky130_fd_sc_hd__o21ai_1 _3347_ (.A1(_1624_),
    .A2(_1651_),
    .B1(_1652_),
    .Y(_0971_));
 sky130_fd_sc_hd__and3_1 _3348_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[10].S.IN1_L2 ),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _3349_ (.A(_1653_),
    .X(_0973_));
 sky130_fd_sc_hd__nand2b_1 _3350_ (.A_N(_0973_),
    .B(_1652_),
    .Y(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3351_ (.A(_1654_),
    .X(_0972_));
 sky130_fd_sc_hd__buf_2 _3352_ (.A(_1582_),
    .X(_1655_));
 sky130_fd_sc_hd__a22oi_4 _3353_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[21].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[21].S.IN1_L3 ),
    .Y(_1656_));
 sky130_fd_sc_hd__and3_1 _3354_ (.A(_1649_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[10].S.IN1_L4 ),
    .X(_1657_));
 sky130_fd_sc_hd__buf_6 _3355_ (.A(_1657_),
    .X(_0975_));
 sky130_fd_sc_hd__o21bai_1 _3356_ (.A1(_1655_),
    .A2(_1656_),
    .B1_N(_0975_),
    .Y(_0974_));
 sky130_fd_sc_hd__a22oi_4 _3357_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[22].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[22].S.IN1_L3 ),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_1 _3358_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[11].S.IN1_L1 ),
    .Y(_1659_));
 sky130_fd_sc_hd__o21ai_1 _3359_ (.A1(_1624_),
    .A2(_1658_),
    .B1(_1659_),
    .Y(_0976_));
 sky130_fd_sc_hd__and3_1 _3360_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[11].S.IN1_L2 ),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3361_ (.A(_1660_),
    .X(_0978_));
 sky130_fd_sc_hd__nand2b_1 _3362_ (.A_N(_0978_),
    .B(_1659_),
    .Y(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _3363_ (.A(_1661_),
    .X(_0977_));
 sky130_fd_sc_hd__a22oi_4 _3364_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[23].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[23].S.IN1_L3 ),
    .Y(_1662_));
 sky130_fd_sc_hd__and3_1 _3365_ (.A(_1649_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[11].S.IN1_L4 ),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(_1663_),
    .X(_0980_));
 sky130_fd_sc_hd__o21bai_1 _3367_ (.A1(_1655_),
    .A2(_1662_),
    .B1_N(_0980_),
    .Y(_0979_));
 sky130_fd_sc_hd__a22oi_4 _3368_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[24].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[24].S.IN1_L3 ),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _3369_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[12].S.IN1_L1 ),
    .Y(_1665_));
 sky130_fd_sc_hd__o21ai_1 _3370_ (.A1(_1624_),
    .A2(_1664_),
    .B1(_1665_),
    .Y(_0981_));
 sky130_fd_sc_hd__and3_1 _3371_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[12].S.IN1_L2 ),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1666_),
    .X(_0983_));
 sky130_fd_sc_hd__nand2b_1 _3373_ (.A_N(_0983_),
    .B(_1665_),
    .Y(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1667_),
    .X(_0982_));
 sky130_fd_sc_hd__a22oi_2 _3375_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[25].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[25].S.IN1_L3 ),
    .Y(_1668_));
 sky130_fd_sc_hd__and3_1 _3376_ (.A(_1649_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[12].S.IN1_L4 ),
    .X(_1669_));
 sky130_fd_sc_hd__buf_6 _3377_ (.A(_1669_),
    .X(_0985_));
 sky130_fd_sc_hd__o21bai_1 _3378_ (.A1(_1655_),
    .A2(_1668_),
    .B1_N(_0985_),
    .Y(_0984_));
 sky130_fd_sc_hd__a22oi_2 _3379_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[26].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[26].S.IN1_L3 ),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _3380_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[13].S.IN1_L1 ),
    .Y(_1671_));
 sky130_fd_sc_hd__o21ai_1 _3381_ (.A1(_1624_),
    .A2(_1670_),
    .B1(_1671_),
    .Y(_0986_));
 sky130_fd_sc_hd__and3_1 _3382_ (.A(_1636_),
    .B(_1606_),
    .C(\stage_gen[3].mux_gen[13].S.IN1_L2 ),
    .X(_1672_));
 sky130_fd_sc_hd__clkbuf_1 _3383_ (.A(_1672_),
    .X(_0988_));
 sky130_fd_sc_hd__nand2b_1 _3384_ (.A_N(_0988_),
    .B(_1671_),
    .Y(_1673_));
 sky130_fd_sc_hd__clkbuf_1 _3385_ (.A(_1673_),
    .X(_0987_));
 sky130_fd_sc_hd__a22oi_1 _3386_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[27].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[27].S.IN1_L3 ),
    .Y(_1674_));
 sky130_fd_sc_hd__and3_1 _3387_ (.A(_1649_),
    .B(_1610_),
    .C(\stage_gen[3].mux_gen[13].S.IN1_L4 ),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3388_ (.A(_1675_),
    .X(_0990_));
 sky130_fd_sc_hd__o21bai_1 _3389_ (.A1(_1655_),
    .A2(_1674_),
    .B1_N(_0990_),
    .Y(_0989_));
 sky130_fd_sc_hd__a22oi_1 _3390_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[28].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[28].S.IN1_L3 ),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _3391_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[14].S.IN1_L1 ),
    .Y(_1677_));
 sky130_fd_sc_hd__o21ai_1 _3392_ (.A1(_1624_),
    .A2(_1676_),
    .B1(_1677_),
    .Y(_0991_));
 sky130_fd_sc_hd__buf_2 _3393_ (.A(_1360_),
    .X(_1678_));
 sky130_fd_sc_hd__and3_1 _3394_ (.A(_1636_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[14].S.IN1_L2 ),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3395_ (.A(_1679_),
    .X(_0993_));
 sky130_fd_sc_hd__nand2b_1 _3396_ (.A_N(_0993_),
    .B(_1677_),
    .Y(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _3397_ (.A(_1680_),
    .X(_0992_));
 sky130_fd_sc_hd__a22oi_2 _3398_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[29].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[29].S.IN1_L3 ),
    .Y(_1681_));
 sky130_fd_sc_hd__buf_6 _3399_ (.A(_1384_),
    .X(_1682_));
 sky130_fd_sc_hd__buf_2 _3400_ (.A(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__and3_1 _3401_ (.A(_1649_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[14].S.IN1_L4 ),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _3402_ (.A(_1684_),
    .X(_0995_));
 sky130_fd_sc_hd__o21bai_1 _3403_ (.A1(_1655_),
    .A2(_1681_),
    .B1_N(_0995_),
    .Y(_0994_));
 sky130_fd_sc_hd__a22oi_1 _3404_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[30].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[30].S.IN1_L3 ),
    .Y(_1685_));
 sky130_fd_sc_hd__nand2_1 _3405_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[15].S.IN1_L1 ),
    .Y(_1686_));
 sky130_fd_sc_hd__o21ai_1 _3406_ (.A1(_1624_),
    .A2(_1685_),
    .B1(_1686_),
    .Y(_0996_));
 sky130_fd_sc_hd__and3_1 _3407_ (.A(_1636_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[15].S.IN1_L2 ),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _3408_ (.A(_1687_),
    .X(_0998_));
 sky130_fd_sc_hd__nand2b_1 _3409_ (.A_N(_0998_),
    .B(_1686_),
    .Y(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1688_),
    .X(_0997_));
 sky130_fd_sc_hd__a22oi_1 _3411_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[31].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[31].S.IN1_L3 ),
    .Y(_1689_));
 sky130_fd_sc_hd__and3_1 _3412_ (.A(_1649_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[15].S.IN1_L4 ),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _3413_ (.A(_1690_),
    .X(_1000_));
 sky130_fd_sc_hd__o21bai_1 _3414_ (.A1(_1655_),
    .A2(_1689_),
    .B1_N(_1000_),
    .Y(_0999_));
 sky130_fd_sc_hd__a22oi_2 _3415_ (.A1(_1625_),
    .A2(\stage_gen[2].mux_gen[32].S.IN1_L5 ),
    .B1(_1626_),
    .B2(\stage_gen[2].mux_gen[32].S.IN1_L3 ),
    .Y(_1691_));
 sky130_fd_sc_hd__nand2_1 _3416_ (.A(_1628_),
    .B(\stage_gen[3].mux_gen[16].S.IN1_L1 ),
    .Y(_1692_));
 sky130_fd_sc_hd__o21ai_1 _3417_ (.A1(_1624_),
    .A2(_1691_),
    .B1(_1692_),
    .Y(_1001_));
 sky130_fd_sc_hd__and3_1 _3418_ (.A(_1636_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[16].S.IN1_L2 ),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _3419_ (.A(_1693_),
    .X(_1003_));
 sky130_fd_sc_hd__nand2b_1 _3420_ (.A_N(_1003_),
    .B(_1692_),
    .Y(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _3421_ (.A(_1694_),
    .X(_1002_));
 sky130_fd_sc_hd__a22oi_1 _3422_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[33].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[33].S.IN1_L3 ),
    .Y(_1695_));
 sky130_fd_sc_hd__and3_1 _3423_ (.A(_1649_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[16].S.IN1_L4 ),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _3424_ (.A(_1696_),
    .X(_1005_));
 sky130_fd_sc_hd__o21bai_1 _3425_ (.A1(_1655_),
    .A2(_1695_),
    .B1_N(_1005_),
    .Y(_1004_));
 sky130_fd_sc_hd__buf_2 _3426_ (.A(_1582_),
    .X(_1697_));
 sky130_fd_sc_hd__buf_4 _3427_ (.A(_1387_),
    .X(_1698_));
 sky130_fd_sc_hd__buf_4 _3428_ (.A(_1569_),
    .X(_1699_));
 sky130_fd_sc_hd__a22oi_2 _3429_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[34].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[34].S.IN1_L3 ),
    .Y(_1700_));
 sky130_fd_sc_hd__buf_2 _3430_ (.A(_1574_),
    .X(_1701_));
 sky130_fd_sc_hd__nand2_1 _3431_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[17].S.IN1_L1 ),
    .Y(_1702_));
 sky130_fd_sc_hd__o21ai_1 _3432_ (.A1(_1697_),
    .A2(_1700_),
    .B1(_1702_),
    .Y(_1006_));
 sky130_fd_sc_hd__and3_1 _3433_ (.A(_1636_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[17].S.IN1_L2 ),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _3434_ (.A(_1703_),
    .X(_1008_));
 sky130_fd_sc_hd__nand2b_1 _3435_ (.A_N(_1008_),
    .B(_1702_),
    .Y(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3436_ (.A(_1704_),
    .X(_1007_));
 sky130_fd_sc_hd__a22oi_1 _3437_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[35].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[35].S.IN1_L3 ),
    .Y(_1705_));
 sky130_fd_sc_hd__and3_1 _3438_ (.A(_1649_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[17].S.IN1_L4 ),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _3439_ (.A(_1706_),
    .X(_1010_));
 sky130_fd_sc_hd__o21bai_1 _3440_ (.A1(_1655_),
    .A2(_1705_),
    .B1_N(_1010_),
    .Y(_1009_));
 sky130_fd_sc_hd__a22oi_2 _3441_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[36].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[36].S.IN1_L3 ),
    .Y(_1707_));
 sky130_fd_sc_hd__nand2_1 _3442_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[18].S.IN1_L1 ),
    .Y(_1708_));
 sky130_fd_sc_hd__o21ai_1 _3443_ (.A1(_1697_),
    .A2(_1707_),
    .B1(_1708_),
    .Y(_1011_));
 sky130_fd_sc_hd__buf_2 _3444_ (.A(_1578_),
    .X(_1709_));
 sky130_fd_sc_hd__and3_1 _3445_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[18].S.IN1_L2 ),
    .X(_1710_));
 sky130_fd_sc_hd__clkbuf_1 _3446_ (.A(_1710_),
    .X(_1013_));
 sky130_fd_sc_hd__nand2b_1 _3447_ (.A_N(_1013_),
    .B(_1708_),
    .Y(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3448_ (.A(_1711_),
    .X(_1012_));
 sky130_fd_sc_hd__a22oi_2 _3449_ (.A1(_1646_),
    .A2(\stage_gen[2].mux_gen[37].S.IN1_L5 ),
    .B1(_1647_),
    .B2(\stage_gen[2].mux_gen[37].S.IN1_L3 ),
    .Y(_1712_));
 sky130_fd_sc_hd__and3_1 _3450_ (.A(_1649_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[18].S.IN1_L4 ),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _3451_ (.A(_1713_),
    .X(_1015_));
 sky130_fd_sc_hd__o21bai_1 _3452_ (.A1(_1655_),
    .A2(_1712_),
    .B1_N(_1015_),
    .Y(_1014_));
 sky130_fd_sc_hd__a22oi_1 _3453_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[38].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[38].S.IN1_L3 ),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2_1 _3454_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[19].S.IN1_L1 ),
    .Y(_1715_));
 sky130_fd_sc_hd__o21ai_1 _3455_ (.A1(_1697_),
    .A2(_1714_),
    .B1(_1715_),
    .Y(_1016_));
 sky130_fd_sc_hd__and3_1 _3456_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[19].S.IN1_L2 ),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3457_ (.A(_1716_),
    .X(_1018_));
 sky130_fd_sc_hd__nand2b_1 _3458_ (.A_N(_1018_),
    .B(_1715_),
    .Y(_1717_));
 sky130_fd_sc_hd__clkbuf_1 _3459_ (.A(_1717_),
    .X(_1017_));
 sky130_fd_sc_hd__buf_4 _3460_ (.A(_1387_),
    .X(_1718_));
 sky130_fd_sc_hd__buf_4 _3461_ (.A(_1570_),
    .X(_1719_));
 sky130_fd_sc_hd__a22oi_1 _3462_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[39].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[39].S.IN1_L3 ),
    .Y(_1720_));
 sky130_fd_sc_hd__clkbuf_2 _3463_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .X(_1721_));
 sky130_fd_sc_hd__and3_1 _3464_ (.A(_1721_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[19].S.IN1_L4 ),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1722_),
    .X(_1020_));
 sky130_fd_sc_hd__o21bai_1 _3466_ (.A1(_1655_),
    .A2(_1720_),
    .B1_N(_1020_),
    .Y(_1019_));
 sky130_fd_sc_hd__a22oi_2 _3467_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[40].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[40].S.IN1_L3 ),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _3468_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[20].S.IN1_L1 ),
    .Y(_1724_));
 sky130_fd_sc_hd__o21ai_1 _3469_ (.A1(_1697_),
    .A2(_1723_),
    .B1(_1724_),
    .Y(_1026_));
 sky130_fd_sc_hd__and3_1 _3470_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[20].S.IN1_L2 ),
    .X(_1725_));
 sky130_fd_sc_hd__clkbuf_1 _3471_ (.A(_1725_),
    .X(_1028_));
 sky130_fd_sc_hd__nand2b_1 _3472_ (.A_N(_1028_),
    .B(_1724_),
    .Y(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _3473_ (.A(_1726_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_4 _3474_ (.A(_1582_),
    .X(_1727_));
 sky130_fd_sc_hd__a22oi_1 _3475_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[41].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[41].S.IN1_L3 ),
    .Y(_1728_));
 sky130_fd_sc_hd__and3_1 _3476_ (.A(_1721_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[20].S.IN1_L4 ),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _3477_ (.A(_1729_),
    .X(_1030_));
 sky130_fd_sc_hd__o21bai_1 _3478_ (.A1(_1727_),
    .A2(_1728_),
    .B1_N(_1030_),
    .Y(_1029_));
 sky130_fd_sc_hd__a22oi_1 _3479_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[42].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[42].S.IN1_L3 ),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[21].S.IN1_L1 ),
    .Y(_1731_));
 sky130_fd_sc_hd__o21ai_1 _3481_ (.A1(_1697_),
    .A2(_1730_),
    .B1(_1731_),
    .Y(_1031_));
 sky130_fd_sc_hd__and3_1 _3482_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[21].S.IN1_L2 ),
    .X(_1732_));
 sky130_fd_sc_hd__clkbuf_1 _3483_ (.A(_1732_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2b_1 _3484_ (.A_N(_1033_),
    .B(_1731_),
    .Y(_1733_));
 sky130_fd_sc_hd__clkbuf_1 _3485_ (.A(_1733_),
    .X(_1032_));
 sky130_fd_sc_hd__a22oi_1 _3486_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[43].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[43].S.IN1_L3 ),
    .Y(_1734_));
 sky130_fd_sc_hd__and3_1 _3487_ (.A(_1721_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[21].S.IN1_L4 ),
    .X(_1735_));
 sky130_fd_sc_hd__clkbuf_1 _3488_ (.A(_1735_),
    .X(_1035_));
 sky130_fd_sc_hd__o21bai_1 _3489_ (.A1(_1727_),
    .A2(_1734_),
    .B1_N(_1035_),
    .Y(_1034_));
 sky130_fd_sc_hd__a22oi_2 _3490_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[44].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[44].S.IN1_L3 ),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _3491_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[22].S.IN1_L1 ),
    .Y(_1737_));
 sky130_fd_sc_hd__o21ai_1 _3492_ (.A1(_1697_),
    .A2(_1736_),
    .B1(_1737_),
    .Y(_1036_));
 sky130_fd_sc_hd__and3_1 _3493_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[22].S.IN1_L2 ),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _3494_ (.A(_1738_),
    .X(_1038_));
 sky130_fd_sc_hd__nand2b_1 _3495_ (.A_N(_1038_),
    .B(_1737_),
    .Y(_1739_));
 sky130_fd_sc_hd__clkbuf_1 _3496_ (.A(_1739_),
    .X(_1037_));
 sky130_fd_sc_hd__a22oi_1 _3497_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[45].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[45].S.IN1_L3 ),
    .Y(_1740_));
 sky130_fd_sc_hd__and3_1 _3498_ (.A(_1721_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[22].S.IN1_L4 ),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1741_),
    .X(_1040_));
 sky130_fd_sc_hd__o21bai_1 _3500_ (.A1(_1727_),
    .A2(_1740_),
    .B1_N(_1040_),
    .Y(_1039_));
 sky130_fd_sc_hd__a22oi_1 _3501_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[46].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[46].S.IN1_L3 ),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _3502_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[23].S.IN1_L1 ),
    .Y(_1743_));
 sky130_fd_sc_hd__o21ai_1 _3503_ (.A1(_1697_),
    .A2(_1742_),
    .B1(_1743_),
    .Y(_1041_));
 sky130_fd_sc_hd__and3_1 _3504_ (.A(_1709_),
    .B(_1678_),
    .C(\stage_gen[3].mux_gen[23].S.IN1_L2 ),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(_1744_),
    .X(_1043_));
 sky130_fd_sc_hd__nand2b_1 _3506_ (.A_N(_1043_),
    .B(_1743_),
    .Y(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _3507_ (.A(_1745_),
    .X(_1042_));
 sky130_fd_sc_hd__a22oi_1 _3508_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[47].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[47].S.IN1_L3 ),
    .Y(_1746_));
 sky130_fd_sc_hd__and3_1 _3509_ (.A(_1721_),
    .B(_1683_),
    .C(\stage_gen[3].mux_gen[23].S.IN1_L4 ),
    .X(_1747_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_1747_),
    .X(_1045_));
 sky130_fd_sc_hd__o21bai_1 _3511_ (.A1(_1727_),
    .A2(_1746_),
    .B1_N(_1045_),
    .Y(_1044_));
 sky130_fd_sc_hd__a22oi_4 _3512_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[48].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[48].S.IN1_L3 ),
    .Y(_1748_));
 sky130_fd_sc_hd__nand2_1 _3513_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[24].S.IN1_L1 ),
    .Y(_1749_));
 sky130_fd_sc_hd__o21ai_1 _3514_ (.A1(_1697_),
    .A2(_1748_),
    .B1(_1749_),
    .Y(_1046_));
 sky130_fd_sc_hd__buf_4 _3515_ (.A(_1360_),
    .X(_1750_));
 sky130_fd_sc_hd__and3_1 _3516_ (.A(_1709_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[24].S.IN1_L2 ),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_1751_),
    .X(_1048_));
 sky130_fd_sc_hd__nand2b_1 _3518_ (.A_N(_1048_),
    .B(_1749_),
    .Y(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(_1752_),
    .X(_1047_));
 sky130_fd_sc_hd__a22oi_2 _3520_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[49].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[49].S.IN1_L3 ),
    .Y(_1753_));
 sky130_fd_sc_hd__buf_4 _3521_ (.A(_1682_),
    .X(_1754_));
 sky130_fd_sc_hd__and3_1 _3522_ (.A(_1721_),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[24].S.IN1_L4 ),
    .X(_1755_));
 sky130_fd_sc_hd__clkbuf_1 _3523_ (.A(_1755_),
    .X(_1050_));
 sky130_fd_sc_hd__o21bai_1 _3524_ (.A1(_1727_),
    .A2(_1753_),
    .B1_N(_1050_),
    .Y(_1049_));
 sky130_fd_sc_hd__a22oi_4 _3525_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[50].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[50].S.IN1_L3 ),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _3526_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[25].S.IN1_L1 ),
    .Y(_1757_));
 sky130_fd_sc_hd__o21ai_1 _3527_ (.A1(_1697_),
    .A2(_1756_),
    .B1(_1757_),
    .Y(_1051_));
 sky130_fd_sc_hd__and3_1 _3528_ (.A(_1709_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[25].S.IN1_L2 ),
    .X(_1758_));
 sky130_fd_sc_hd__clkbuf_1 _3529_ (.A(_1758_),
    .X(_1053_));
 sky130_fd_sc_hd__nand2b_1 _3530_ (.A_N(_1053_),
    .B(_1757_),
    .Y(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _3531_ (.A(_1759_),
    .X(_1052_));
 sky130_fd_sc_hd__a22oi_2 _3532_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[51].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[51].S.IN1_L3 ),
    .Y(_1760_));
 sky130_fd_sc_hd__and3_1 _3533_ (.A(_1721_),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[25].S.IN1_L4 ),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _3534_ (.A(_1761_),
    .X(_1055_));
 sky130_fd_sc_hd__o21bai_1 _3535_ (.A1(_1727_),
    .A2(_1760_),
    .B1_N(_1055_),
    .Y(_1054_));
 sky130_fd_sc_hd__a22oi_2 _3536_ (.A1(_1698_),
    .A2(\stage_gen[2].mux_gen[52].S.IN1_L5 ),
    .B1(_1699_),
    .B2(\stage_gen[2].mux_gen[52].S.IN1_L3 ),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _3537_ (.A(_1701_),
    .B(\stage_gen[3].mux_gen[26].S.IN1_L1 ),
    .Y(_1763_));
 sky130_fd_sc_hd__o21ai_1 _3538_ (.A1(_1697_),
    .A2(_1762_),
    .B1(_1763_),
    .Y(_1056_));
 sky130_fd_sc_hd__and3_1 _3539_ (.A(_1709_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[26].S.IN1_L2 ),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_1764_),
    .X(_1058_));
 sky130_fd_sc_hd__nand2b_1 _3541_ (.A_N(_1058_),
    .B(_1763_),
    .Y(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _3542_ (.A(_1765_),
    .X(_1057_));
 sky130_fd_sc_hd__a22oi_2 _3543_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[53].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[53].S.IN1_L3 ),
    .Y(_1766_));
 sky130_fd_sc_hd__and3_1 _3544_ (.A(_1721_),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[26].S.IN1_L4 ),
    .X(_1767_));
 sky130_fd_sc_hd__clkbuf_1 _3545_ (.A(_1767_),
    .X(_1060_));
 sky130_fd_sc_hd__o21bai_1 _3546_ (.A1(_1727_),
    .A2(_1766_),
    .B1_N(_1060_),
    .Y(_1059_));
 sky130_fd_sc_hd__a22oi_2 _3547_ (.A1(_1388_),
    .A2(\stage_gen[2].mux_gen[54].S.IN1_L5 ),
    .B1(_1570_),
    .B2(\stage_gen[2].mux_gen[54].S.IN1_L3 ),
    .Y(_1768_));
 sky130_fd_sc_hd__nand2_1 _3548_ (.A(_1575_),
    .B(\stage_gen[3].mux_gen[27].S.IN1_L1 ),
    .Y(_1769_));
 sky130_fd_sc_hd__o21ai_1 _3549_ (.A1(_1582_),
    .A2(_1768_),
    .B1(_1769_),
    .Y(_1061_));
 sky130_fd_sc_hd__and3_1 _3550_ (.A(_1709_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[27].S.IN1_L2 ),
    .X(_1770_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1770_),
    .X(_1063_));
 sky130_fd_sc_hd__nand2b_1 _3552_ (.A_N(_1063_),
    .B(_1769_),
    .Y(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1771_),
    .X(_1062_));
 sky130_fd_sc_hd__a22oi_2 _3554_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[55].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[55].S.IN1_L3 ),
    .Y(_1772_));
 sky130_fd_sc_hd__and3_1 _3555_ (.A(_1721_),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[27].S.IN1_L4 ),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _3556_ (.A(_1773_),
    .X(_1065_));
 sky130_fd_sc_hd__o21bai_1 _3557_ (.A1(_1727_),
    .A2(_1772_),
    .B1_N(_1065_),
    .Y(_1064_));
 sky130_fd_sc_hd__a22oi_2 _3558_ (.A1(_1388_),
    .A2(\stage_gen[2].mux_gen[56].S.IN1_L5 ),
    .B1(_1570_),
    .B2(\stage_gen[2].mux_gen[56].S.IN1_L3 ),
    .Y(_1774_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(_1575_),
    .B(\stage_gen[3].mux_gen[28].S.IN1_L1 ),
    .Y(_1775_));
 sky130_fd_sc_hd__o21ai_1 _3560_ (.A1(_1582_),
    .A2(_1774_),
    .B1(_1775_),
    .Y(_1066_));
 sky130_fd_sc_hd__and3_1 _3561_ (.A(_1578_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[28].S.IN1_L2 ),
    .X(_1776_));
 sky130_fd_sc_hd__clkbuf_1 _3562_ (.A(_1776_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2b_1 _3563_ (.A_N(_1068_),
    .B(_1775_),
    .Y(_1777_));
 sky130_fd_sc_hd__clkbuf_1 _3564_ (.A(_1777_),
    .X(_1067_));
 sky130_fd_sc_hd__a22oi_2 _3565_ (.A1(_1718_),
    .A2(\stage_gen[2].mux_gen[57].S.IN1_L5 ),
    .B1(_1719_),
    .B2(\stage_gen[2].mux_gen[57].S.IN1_L3 ),
    .Y(_1778_));
 sky130_fd_sc_hd__and3_1 _3566_ (.A(_1721_),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[28].S.IN1_L4 ),
    .X(_1779_));
 sky130_fd_sc_hd__clkbuf_1 _3567_ (.A(_1779_),
    .X(_1070_));
 sky130_fd_sc_hd__o21bai_1 _3568_ (.A1(_1727_),
    .A2(_1778_),
    .B1_N(_1070_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22oi_2 _3569_ (.A1(_1388_),
    .A2(\stage_gen[2].mux_gen[58].S.IN1_L5 ),
    .B1(_1570_),
    .B2(\stage_gen[2].mux_gen[58].S.IN1_L3 ),
    .Y(_1780_));
 sky130_fd_sc_hd__nand2_1 _3570_ (.A(_1575_),
    .B(\stage_gen[3].mux_gen[29].S.IN1_L1 ),
    .Y(_1781_));
 sky130_fd_sc_hd__o21ai_1 _3571_ (.A1(_1582_),
    .A2(_1780_),
    .B1(_1781_),
    .Y(_1071_));
 sky130_fd_sc_hd__and3_1 _3572_ (.A(_1578_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[29].S.IN1_L2 ),
    .X(_1782_));
 sky130_fd_sc_hd__clkbuf_1 _3573_ (.A(_1782_),
    .X(_1073_));
 sky130_fd_sc_hd__nand2b_1 _3574_ (.A_N(_1073_),
    .B(_1781_),
    .Y(_1783_));
 sky130_fd_sc_hd__clkbuf_1 _3575_ (.A(_1783_),
    .X(_1072_));
 sky130_fd_sc_hd__a22oi_4 _3576_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[59].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[59].S.IN1_L3 ),
    .Y(_1784_));
 sky130_fd_sc_hd__and3_1 _3577_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[29].S.IN1_L4 ),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _3578_ (.A(_1785_),
    .X(_1075_));
 sky130_fd_sc_hd__o21bai_1 _3579_ (.A1(_1727_),
    .A2(_1784_),
    .B1_N(_1075_),
    .Y(_1074_));
 sky130_fd_sc_hd__a22oi_2 _3580_ (.A1(_1388_),
    .A2(\stage_gen[2].mux_gen[60].S.IN1_L5 ),
    .B1(_1570_),
    .B2(\stage_gen[2].mux_gen[60].S.IN1_L3 ),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(_1575_),
    .B(\stage_gen[3].mux_gen[30].S.IN1_L1 ),
    .Y(_1787_));
 sky130_fd_sc_hd__o21ai_1 _3582_ (.A1(_1582_),
    .A2(_1786_),
    .B1(_1787_),
    .Y(_1081_));
 sky130_fd_sc_hd__and3_1 _3583_ (.A(_1578_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[30].S.IN1_L2 ),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3584_ (.A(_1788_),
    .X(_1083_));
 sky130_fd_sc_hd__nand2b_1 _3585_ (.A_N(_1083_),
    .B(_1787_),
    .Y(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _3586_ (.A(_1789_),
    .X(_1082_));
 sky130_fd_sc_hd__a22oi_2 _3587_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[61].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[61].S.IN1_L3 ),
    .Y(_1790_));
 sky130_fd_sc_hd__and3_1 _3588_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[30].S.IN1_L4 ),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_1 _3589_ (.A(_1791_),
    .X(_1085_));
 sky130_fd_sc_hd__o21bai_1 _3590_ (.A1(_1566_),
    .A2(_1790_),
    .B1_N(_1085_),
    .Y(_1084_));
 sky130_fd_sc_hd__a22oi_2 _3591_ (.A1(_1388_),
    .A2(\stage_gen[2].mux_gen[62].S.IN1_L5 ),
    .B1(_1570_),
    .B2(\stage_gen[2].mux_gen[62].S.IN1_L3 ),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _3592_ (.A(_1575_),
    .B(\stage_gen[3].mux_gen[31].S.IN1_L1 ),
    .Y(_1793_));
 sky130_fd_sc_hd__o21ai_1 _3593_ (.A1(_1582_),
    .A2(_1792_),
    .B1(_1793_),
    .Y(_1086_));
 sky130_fd_sc_hd__and3_1 _3594_ (.A(_1578_),
    .B(_1750_),
    .C(\stage_gen[3].mux_gen[31].S.IN1_L2 ),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _3595_ (.A(_1794_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2b_1 _3596_ (.A_N(_1088_),
    .B(_1793_),
    .Y(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3597_ (.A(_1795_),
    .X(_1087_));
 sky130_fd_sc_hd__a22oi_4 _3598_ (.A1(_1567_),
    .A2(\stage_gen[2].mux_gen[63].S.IN1_L5 ),
    .B1(_1571_),
    .B2(\stage_gen[2].mux_gen[63].S.IN1_L3 ),
    .Y(_1796_));
 sky130_fd_sc_hd__and3_1 _3599_ (.A(\stage_gen[3].genblk1.clks.clk_o ),
    .B(_1754_),
    .C(\stage_gen[3].mux_gen[31].S.IN1_L4 ),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _3600_ (.A(_1797_),
    .X(_1090_));
 sky130_fd_sc_hd__o21bai_1 _3601_ (.A1(_1566_),
    .A2(_1796_),
    .B1_N(_1090_),
    .Y(_1089_));
 sky130_fd_sc_hd__clkbuf_2 _3602_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_4 _3603_ (.A(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__buf_4 _3604_ (.A(_1575_),
    .X(_1800_));
 sky130_fd_sc_hd__buf_6 _3605_ (.A(_1360_),
    .X(_1801_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_1579_),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__clkinv_4 _3607_ (.A(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__buf_6 _3608_ (.A(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__a22oi_1 _3609_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[0].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[0].S.IN1_L3 ),
    .Y(_1805_));
 sky130_fd_sc_hd__nand2_1 _3610_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .B(_1682_),
    .Y(_1806_));
 sky130_fd_sc_hd__clkinv_4 _3611_ (.A(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__buf_4 _3612_ (.A(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nand2_1 _3613_ (.A(_1808_),
    .B(\stage_gen[4].mux_gen[0].S.IN1_L1 ),
    .Y(_1809_));
 sky130_fd_sc_hd__o21ai_1 _3614_ (.A1(_1799_),
    .A2(_1805_),
    .B1(_1809_),
    .Y(_1126_));
 sky130_fd_sc_hd__clkinv_2 _3615_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .Y(_1810_));
 sky130_fd_sc_hd__clkbuf_4 _3616_ (.A(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__and3_1 _3617_ (.A(_1811_),
    .B(_1750_),
    .C(\stage_gen[4].mux_gen[0].S.IN1_L2 ),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_1 _3618_ (.A(_1812_),
    .X(_1128_));
 sky130_fd_sc_hd__nand2b_1 _3619_ (.A_N(_1128_),
    .B(_1809_),
    .Y(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3620_ (.A(_1813_),
    .X(_1127_));
 sky130_fd_sc_hd__buf_2 _3621_ (.A(_1798_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _3622_ (.A(_1575_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _3623_ (.A(_1803_),
    .X(_0970_));
 sky130_fd_sc_hd__a22oi_2 _3624_ (.A1(net395),
    .A2(\stage_gen[3].mux_gen[1].S.IN1_L5 ),
    .B1(net299),
    .B2(\stage_gen[3].mux_gen[1].S.IN1_L3 ),
    .Y(_1815_));
 sky130_fd_sc_hd__and3_1 _3625_ (.A(_1798_),
    .B(_1754_),
    .C(\stage_gen[4].mux_gen[0].S.IN1_L4 ),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _3626_ (.A(_1816_),
    .X(_1130_));
 sky130_fd_sc_hd__o21bai_1 _3627_ (.A1(_1814_),
    .A2(_1815_),
    .B1_N(_1130_),
    .Y(_1129_));
 sky130_fd_sc_hd__a22oi_2 _3628_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[2].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[2].S.IN1_L3 ),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(_1808_),
    .B(\stage_gen[4].mux_gen[1].S.IN1_L1 ),
    .Y(_1818_));
 sky130_fd_sc_hd__o21ai_1 _3630_ (.A1(_1799_),
    .A2(_1817_),
    .B1(_1818_),
    .Y(_1163_));
 sky130_fd_sc_hd__and3_1 _3631_ (.A(_1811_),
    .B(_1750_),
    .C(\stage_gen[4].mux_gen[1].S.IN1_L2 ),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _3632_ (.A(_1819_),
    .X(_1165_));
 sky130_fd_sc_hd__nand2b_1 _3633_ (.A_N(_1165_),
    .B(_1818_),
    .Y(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _3634_ (.A(_1820_),
    .X(_1164_));
 sky130_fd_sc_hd__a22oi_2 _3635_ (.A1(net394),
    .A2(\stage_gen[3].mux_gen[3].S.IN1_L5 ),
    .B1(net299),
    .B2(\stage_gen[3].mux_gen[3].S.IN1_L3 ),
    .Y(_1821_));
 sky130_fd_sc_hd__and3_1 _3636_ (.A(_1798_),
    .B(_1754_),
    .C(\stage_gen[4].mux_gen[1].S.IN1_L4 ),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _3637_ (.A(_1822_),
    .X(_1167_));
 sky130_fd_sc_hd__o21bai_1 _3638_ (.A1(_1814_),
    .A2(_1821_),
    .B1_N(_1167_),
    .Y(_1166_));
 sky130_fd_sc_hd__a22oi_2 _3639_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[4].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[4].S.IN1_L3 ),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _3640_ (.A(_1808_),
    .B(\stage_gen[4].mux_gen[2].S.IN1_L1 ),
    .Y(_1824_));
 sky130_fd_sc_hd__o21ai_1 _3641_ (.A1(_1799_),
    .A2(_1823_),
    .B1(_1824_),
    .Y(_1168_));
 sky130_fd_sc_hd__buf_2 _3642_ (.A(_1384_),
    .X(_1825_));
 sky130_fd_sc_hd__and3_1 _3643_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[2].S.IN1_L2 ),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _3644_ (.A(_1826_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2b_1 _3645_ (.A_N(_1170_),
    .B(_1824_),
    .Y(_1827_));
 sky130_fd_sc_hd__clkbuf_1 _3646_ (.A(_1827_),
    .X(_1169_));
 sky130_fd_sc_hd__a22oi_2 _3647_ (.A1(net396),
    .A2(\stage_gen[3].mux_gen[5].S.IN1_L5 ),
    .B1(net301),
    .B2(\stage_gen[3].mux_gen[5].S.IN1_L3 ),
    .Y(_1828_));
 sky130_fd_sc_hd__buf_4 _3648_ (.A(_1682_),
    .X(_1829_));
 sky130_fd_sc_hd__and3_1 _3649_ (.A(_1798_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[2].S.IN1_L4 ),
    .X(_1830_));
 sky130_fd_sc_hd__clkbuf_1 _3650_ (.A(_1830_),
    .X(_1172_));
 sky130_fd_sc_hd__o21bai_1 _3651_ (.A1(_1814_),
    .A2(_1828_),
    .B1_N(_1172_),
    .Y(_1171_));
 sky130_fd_sc_hd__buf_2 _3652_ (.A(_1798_),
    .X(_1831_));
 sky130_fd_sc_hd__buf_4 _3653_ (.A(_1575_),
    .X(_1832_));
 sky130_fd_sc_hd__buf_6 _3654_ (.A(_1803_),
    .X(_1833_));
 sky130_fd_sc_hd__a22oi_1 _3655_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[6].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[6].S.IN1_L3 ),
    .Y(_1834_));
 sky130_fd_sc_hd__buf_4 _3656_ (.A(_1807_),
    .X(_1835_));
 sky130_fd_sc_hd__nand2_1 _3657_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[3].S.IN1_L1 ),
    .Y(_1836_));
 sky130_fd_sc_hd__o21ai_1 _3658_ (.A1(_1831_),
    .A2(_1834_),
    .B1(_1836_),
    .Y(_1173_));
 sky130_fd_sc_hd__and3_1 _3659_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[3].S.IN1_L2 ),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _3660_ (.A(_1837_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2b_1 _3661_ (.A_N(_1175_),
    .B(_1836_),
    .Y(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _3662_ (.A(_1838_),
    .X(_1174_));
 sky130_fd_sc_hd__a22oi_1 _3663_ (.A1(net401),
    .A2(\stage_gen[3].mux_gen[7].S.IN1_L5 ),
    .B1(net302),
    .B2(\stage_gen[3].mux_gen[7].S.IN1_L3 ),
    .Y(_1839_));
 sky130_fd_sc_hd__and3_1 _3664_ (.A(_1798_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[3].S.IN1_L4 ),
    .X(_1840_));
 sky130_fd_sc_hd__clkbuf_1 _3665_ (.A(_1840_),
    .X(_1177_));
 sky130_fd_sc_hd__o21bai_1 _3666_ (.A1(_1814_),
    .A2(_1839_),
    .B1_N(_1177_),
    .Y(_1176_));
 sky130_fd_sc_hd__a22oi_1 _3667_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[8].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[8].S.IN1_L3 ),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _3668_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[4].S.IN1_L1 ),
    .Y(_1842_));
 sky130_fd_sc_hd__o21ai_1 _3669_ (.A1(_1831_),
    .A2(_1841_),
    .B1(_1842_),
    .Y(_1178_));
 sky130_fd_sc_hd__and3_1 _3670_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[4].S.IN1_L2 ),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _3671_ (.A(_1843_),
    .X(_1180_));
 sky130_fd_sc_hd__nand2b_1 _3672_ (.A_N(_1180_),
    .B(_1842_),
    .Y(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _3673_ (.A(_1844_),
    .X(_1179_));
 sky130_fd_sc_hd__a22oi_2 _3674_ (.A1(net390),
    .A2(\stage_gen[3].mux_gen[9].S.IN1_L5 ),
    .B1(net296),
    .B2(\stage_gen[3].mux_gen[9].S.IN1_L3 ),
    .Y(_1845_));
 sky130_fd_sc_hd__buf_2 _3675_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .X(_1846_));
 sky130_fd_sc_hd__and3_1 _3676_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[4].S.IN1_L4 ),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _3677_ (.A(_1847_),
    .X(_1182_));
 sky130_fd_sc_hd__o21bai_1 _3678_ (.A1(_1814_),
    .A2(_1845_),
    .B1_N(_1182_),
    .Y(_1181_));
 sky130_fd_sc_hd__a22oi_2 _3679_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[10].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[10].S.IN1_L3 ),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[5].S.IN1_L1 ),
    .Y(_1849_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(_1831_),
    .A2(_1848_),
    .B1(_1849_),
    .Y(_1183_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[5].S.IN1_L2 ),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _3683_ (.A(_1850_),
    .X(_1185_));
 sky130_fd_sc_hd__nand2b_1 _3684_ (.A_N(_1185_),
    .B(_1849_),
    .Y(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _3685_ (.A(_1851_),
    .X(_1184_));
 sky130_fd_sc_hd__a22oi_2 _3686_ (.A1(net389),
    .A2(\stage_gen[3].mux_gen[11].S.IN1_L5 ),
    .B1(net295),
    .B2(\stage_gen[3].mux_gen[11].S.IN1_L3 ),
    .Y(_1852_));
 sky130_fd_sc_hd__and3_1 _3687_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[5].S.IN1_L4 ),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _3688_ (.A(_1853_),
    .X(_1187_));
 sky130_fd_sc_hd__o21bai_1 _3689_ (.A1(_1814_),
    .A2(_1852_),
    .B1_N(_1187_),
    .Y(_1186_));
 sky130_fd_sc_hd__a22oi_2 _3690_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[12].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[12].S.IN1_L3 ),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[6].S.IN1_L1 ),
    .Y(_1855_));
 sky130_fd_sc_hd__o21ai_1 _3692_ (.A1(_1831_),
    .A2(_1854_),
    .B1(_1855_),
    .Y(_1188_));
 sky130_fd_sc_hd__and3_1 _3693_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[6].S.IN1_L2 ),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _3694_ (.A(_1856_),
    .X(_1190_));
 sky130_fd_sc_hd__nand2b_1 _3695_ (.A_N(_1190_),
    .B(_1855_),
    .Y(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _3696_ (.A(_1857_),
    .X(_1189_));
 sky130_fd_sc_hd__a22oi_4 _3697_ (.A1(net389),
    .A2(\stage_gen[3].mux_gen[13].S.IN1_L5 ),
    .B1(net295),
    .B2(\stage_gen[3].mux_gen[13].S.IN1_L3 ),
    .Y(_1858_));
 sky130_fd_sc_hd__and3_1 _3698_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[6].S.IN1_L4 ),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _3699_ (.A(_1859_),
    .X(_1192_));
 sky130_fd_sc_hd__o21bai_1 _3700_ (.A1(_1814_),
    .A2(_1858_),
    .B1_N(_1192_),
    .Y(_1191_));
 sky130_fd_sc_hd__a22oi_2 _3701_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[14].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[14].S.IN1_L3 ),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _3702_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[7].S.IN1_L1 ),
    .Y(_1861_));
 sky130_fd_sc_hd__o21ai_1 _3703_ (.A1(_1831_),
    .A2(_1860_),
    .B1(_1861_),
    .Y(_1193_));
 sky130_fd_sc_hd__and3_1 _3704_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[7].S.IN1_L2 ),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _3705_ (.A(_1862_),
    .X(_1195_));
 sky130_fd_sc_hd__nand2b_1 _3706_ (.A_N(_1195_),
    .B(_1861_),
    .Y(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _3707_ (.A(_1863_),
    .X(_1194_));
 sky130_fd_sc_hd__a22oi_2 _3708_ (.A1(net390),
    .A2(\stage_gen[3].mux_gen[15].S.IN1_L5 ),
    .B1(net296),
    .B2(\stage_gen[3].mux_gen[15].S.IN1_L3 ),
    .Y(_1864_));
 sky130_fd_sc_hd__and3_1 _3709_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[7].S.IN1_L4 ),
    .X(_1865_));
 sky130_fd_sc_hd__clkbuf_1 _3710_ (.A(_1865_),
    .X(_1197_));
 sky130_fd_sc_hd__o21bai_1 _3711_ (.A1(_1814_),
    .A2(_1864_),
    .B1_N(_1197_),
    .Y(_1196_));
 sky130_fd_sc_hd__a22oi_1 _3712_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[16].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[16].S.IN1_L3 ),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _3713_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[8].S.IN1_L1 ),
    .Y(_1867_));
 sky130_fd_sc_hd__o21ai_1 _3714_ (.A1(_1831_),
    .A2(_1866_),
    .B1(_1867_),
    .Y(_1198_));
 sky130_fd_sc_hd__and3_1 _3715_ (.A(_1811_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[8].S.IN1_L2 ),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _3716_ (.A(_1868_),
    .X(_1200_));
 sky130_fd_sc_hd__nand2b_1 _3717_ (.A_N(_1200_),
    .B(_1867_),
    .Y(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _3718_ (.A(_1869_),
    .X(_1199_));
 sky130_fd_sc_hd__a22oi_2 _3719_ (.A1(net391),
    .A2(\stage_gen[3].mux_gen[17].S.IN1_L5 ),
    .B1(net297),
    .B2(\stage_gen[3].mux_gen[17].S.IN1_L3 ),
    .Y(_1870_));
 sky130_fd_sc_hd__and3_1 _3720_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[8].S.IN1_L4 ),
    .X(_1871_));
 sky130_fd_sc_hd__clkbuf_1 _3721_ (.A(_1871_),
    .X(_1202_));
 sky130_fd_sc_hd__o21bai_1 _3722_ (.A1(_1814_),
    .A2(_1870_),
    .B1_N(_1202_),
    .Y(_1201_));
 sky130_fd_sc_hd__a22oi_1 _3723_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[18].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[18].S.IN1_L3 ),
    .Y(_1872_));
 sky130_fd_sc_hd__nand2_1 _3724_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[9].S.IN1_L1 ),
    .Y(_1873_));
 sky130_fd_sc_hd__o21ai_1 _3725_ (.A1(_1831_),
    .A2(_1872_),
    .B1(_1873_),
    .Y(_1203_));
 sky130_fd_sc_hd__and3_1 _3726_ (.A(_1810_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[9].S.IN1_L2 ),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _3727_ (.A(_1874_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2b_1 _3728_ (.A_N(_1205_),
    .B(_1873_),
    .Y(_1875_));
 sky130_fd_sc_hd__clkbuf_1 _3729_ (.A(_1875_),
    .X(_1204_));
 sky130_fd_sc_hd__a22oi_1 _3730_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[19].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[19].S.IN1_L3 ),
    .Y(_1876_));
 sky130_fd_sc_hd__and3_1 _3731_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[9].S.IN1_L4 ),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _3732_ (.A(_1877_),
    .X(_1207_));
 sky130_fd_sc_hd__o21bai_1 _3733_ (.A1(_1814_),
    .A2(_1876_),
    .B1_N(_1207_),
    .Y(_1206_));
 sky130_fd_sc_hd__a22oi_1 _3734_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[20].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[20].S.IN1_L3 ),
    .Y(_1878_));
 sky130_fd_sc_hd__nand2_1 _3735_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[10].S.IN1_L1 ),
    .Y(_1879_));
 sky130_fd_sc_hd__o21ai_1 _3736_ (.A1(_1831_),
    .A2(_1878_),
    .B1(_1879_),
    .Y(_1133_));
 sky130_fd_sc_hd__and3_1 _3737_ (.A(_1810_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[10].S.IN1_L2 ),
    .X(_1880_));
 sky130_fd_sc_hd__clkbuf_1 _3738_ (.A(_1880_),
    .X(_1135_));
 sky130_fd_sc_hd__nand2b_1 _3739_ (.A_N(_1135_),
    .B(_1879_),
    .Y(_1881_));
 sky130_fd_sc_hd__clkbuf_1 _3740_ (.A(_1881_),
    .X(_1134_));
 sky130_fd_sc_hd__a22oi_1 _3741_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[21].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[21].S.IN1_L3 ),
    .Y(_1882_));
 sky130_fd_sc_hd__and3_1 _3742_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[10].S.IN1_L4 ),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _3743_ (.A(_1883_),
    .X(_1137_));
 sky130_fd_sc_hd__o21bai_1 _3744_ (.A1(_1799_),
    .A2(_1882_),
    .B1_N(_1137_),
    .Y(_1136_));
 sky130_fd_sc_hd__a22oi_1 _3745_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[22].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[22].S.IN1_L3 ),
    .Y(_1884_));
 sky130_fd_sc_hd__nand2_1 _3746_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[11].S.IN1_L1 ),
    .Y(_1885_));
 sky130_fd_sc_hd__o21ai_1 _3747_ (.A1(_1831_),
    .A2(_1884_),
    .B1(_1885_),
    .Y(_1138_));
 sky130_fd_sc_hd__and3_1 _3748_ (.A(_1810_),
    .B(_1825_),
    .C(\stage_gen[4].mux_gen[11].S.IN1_L2 ),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _3749_ (.A(_1886_),
    .X(_1140_));
 sky130_fd_sc_hd__nand2b_1 _3750_ (.A_N(_1140_),
    .B(_1885_),
    .Y(_1887_));
 sky130_fd_sc_hd__clkbuf_1 _3751_ (.A(_1887_),
    .X(_1139_));
 sky130_fd_sc_hd__a22oi_1 _3752_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[23].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[23].S.IN1_L3 ),
    .Y(_1888_));
 sky130_fd_sc_hd__and3_1 _3753_ (.A(_1846_),
    .B(_1829_),
    .C(\stage_gen[4].mux_gen[11].S.IN1_L4 ),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _3754_ (.A(_1889_),
    .X(_1142_));
 sky130_fd_sc_hd__o21bai_1 _3755_ (.A1(_1799_),
    .A2(_1888_),
    .B1_N(_1142_),
    .Y(_1141_));
 sky130_fd_sc_hd__a22oi_1 _3756_ (.A1(_1832_),
    .A2(\stage_gen[3].mux_gen[24].S.IN1_L5 ),
    .B1(_1833_),
    .B2(\stage_gen[3].mux_gen[24].S.IN1_L3 ),
    .Y(_1890_));
 sky130_fd_sc_hd__nand2_1 _3757_ (.A(_1835_),
    .B(\stage_gen[4].mux_gen[12].S.IN1_L1 ),
    .Y(_1891_));
 sky130_fd_sc_hd__o21ai_1 _3758_ (.A1(_1831_),
    .A2(_1890_),
    .B1(_1891_),
    .Y(_1143_));
 sky130_fd_sc_hd__buf_4 _3759_ (.A(_1384_),
    .X(_1892_));
 sky130_fd_sc_hd__and3_1 _3760_ (.A(_1810_),
    .B(_1892_),
    .C(\stage_gen[4].mux_gen[12].S.IN1_L2 ),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _3761_ (.A(_1893_),
    .X(_1145_));
 sky130_fd_sc_hd__nand2b_1 _3762_ (.A_N(_1145_),
    .B(_1891_),
    .Y(_1894_));
 sky130_fd_sc_hd__clkbuf_1 _3763_ (.A(_1894_),
    .X(_1144_));
 sky130_fd_sc_hd__a22oi_1 _3764_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[25].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[25].S.IN1_L3 ),
    .Y(_1895_));
 sky130_fd_sc_hd__buf_4 _3765_ (.A(_1682_),
    .X(_1896_));
 sky130_fd_sc_hd__and3_1 _3766_ (.A(_1846_),
    .B(_1896_),
    .C(\stage_gen[4].mux_gen[12].S.IN1_L4 ),
    .X(_1897_));
 sky130_fd_sc_hd__clkbuf_1 _3767_ (.A(_1897_),
    .X(_1147_));
 sky130_fd_sc_hd__o21bai_1 _3768_ (.A1(_1799_),
    .A2(_1895_),
    .B1_N(_1147_),
    .Y(_1146_));
 sky130_fd_sc_hd__a22oi_1 _3769_ (.A1(_1576_),
    .A2(\stage_gen[3].mux_gen[26].S.IN1_L5 ),
    .B1(_1803_),
    .B2(\stage_gen[3].mux_gen[26].S.IN1_L3 ),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _3770_ (.A(_1807_),
    .B(\stage_gen[4].mux_gen[13].S.IN1_L1 ),
    .Y(_1899_));
 sky130_fd_sc_hd__o21ai_1 _3771_ (.A1(_1798_),
    .A2(_1898_),
    .B1(_1899_),
    .Y(_1148_));
 sky130_fd_sc_hd__and3_1 _3772_ (.A(_1810_),
    .B(_1892_),
    .C(\stage_gen[4].mux_gen[13].S.IN1_L2 ),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _3773_ (.A(_1900_),
    .X(_1150_));
 sky130_fd_sc_hd__nand2b_1 _3774_ (.A_N(_1150_),
    .B(_1899_),
    .Y(_1901_));
 sky130_fd_sc_hd__clkbuf_1 _3775_ (.A(_1901_),
    .X(_1149_));
 sky130_fd_sc_hd__a22oi_1 _3776_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[27].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[27].S.IN1_L3 ),
    .Y(_1902_));
 sky130_fd_sc_hd__and3_1 _3777_ (.A(_1846_),
    .B(_1896_),
    .C(\stage_gen[4].mux_gen[13].S.IN1_L4 ),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _3778_ (.A(_1903_),
    .X(_1152_));
 sky130_fd_sc_hd__o21bai_1 _3779_ (.A1(_1799_),
    .A2(_1902_),
    .B1_N(_1152_),
    .Y(_1151_));
 sky130_fd_sc_hd__a22oi_1 _3780_ (.A1(_1576_),
    .A2(\stage_gen[3].mux_gen[28].S.IN1_L5 ),
    .B1(_1803_),
    .B2(\stage_gen[3].mux_gen[28].S.IN1_L3 ),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2_1 _3781_ (.A(_1807_),
    .B(\stage_gen[4].mux_gen[14].S.IN1_L1 ),
    .Y(_1905_));
 sky130_fd_sc_hd__o21ai_1 _3782_ (.A1(_1798_),
    .A2(_1904_),
    .B1(_1905_),
    .Y(_1153_));
 sky130_fd_sc_hd__and3_1 _3783_ (.A(_1810_),
    .B(_1892_),
    .C(\stage_gen[4].mux_gen[14].S.IN1_L2 ),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _3784_ (.A(_1906_),
    .X(_1155_));
 sky130_fd_sc_hd__nand2b_1 _3785_ (.A_N(_1155_),
    .B(_1905_),
    .Y(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _3786_ (.A(_1907_),
    .X(_1154_));
 sky130_fd_sc_hd__a22oi_1 _3787_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[29].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[29].S.IN1_L3 ),
    .Y(_1908_));
 sky130_fd_sc_hd__and3_1 _3788_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[4].mux_gen[14].S.IN1_L4 ),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _3789_ (.A(_1909_),
    .X(_1157_));
 sky130_fd_sc_hd__o21bai_1 _3790_ (.A1(_1799_),
    .A2(_1908_),
    .B1_N(_1157_),
    .Y(_1156_));
 sky130_fd_sc_hd__a22oi_1 _3791_ (.A1(_1576_),
    .A2(\stage_gen[3].mux_gen[30].S.IN1_L5 ),
    .B1(_1803_),
    .B2(\stage_gen[3].mux_gen[30].S.IN1_L3 ),
    .Y(_1910_));
 sky130_fd_sc_hd__nand2_1 _3792_ (.A(_1807_),
    .B(\stage_gen[4].mux_gen[15].S.IN1_L1 ),
    .Y(_1911_));
 sky130_fd_sc_hd__o21ai_1 _3793_ (.A1(_1798_),
    .A2(_1910_),
    .B1(_1911_),
    .Y(_1158_));
 sky130_fd_sc_hd__and3_1 _3794_ (.A(_1810_),
    .B(_1892_),
    .C(\stage_gen[4].mux_gen[15].S.IN1_L2 ),
    .X(_1912_));
 sky130_fd_sc_hd__clkbuf_1 _3795_ (.A(_1912_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2b_1 _3796_ (.A_N(_1160_),
    .B(_1911_),
    .Y(_1913_));
 sky130_fd_sc_hd__clkbuf_1 _3797_ (.A(_1913_),
    .X(_1159_));
 sky130_fd_sc_hd__a22oi_1 _3798_ (.A1(_1800_),
    .A2(\stage_gen[3].mux_gen[31].S.IN1_L5 ),
    .B1(_1804_),
    .B2(\stage_gen[3].mux_gen[31].S.IN1_L3 ),
    .Y(_1914_));
 sky130_fd_sc_hd__and3_1 _3799_ (.A(\stage_gen[4].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[4].mux_gen[15].S.IN1_L4 ),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _3800_ (.A(_1915_),
    .X(_1162_));
 sky130_fd_sc_hd__o21bai_1 _3801_ (.A1(_1799_),
    .A2(_1914_),
    .B1_N(_1162_),
    .Y(_1161_));
 sky130_fd_sc_hd__buf_4 _3802_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .X(_1916_));
 sky130_fd_sc_hd__buf_4 _3803_ (.A(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__clkbuf_1 _3804_ (.A(_1807_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _3805_ (.A(_1810_),
    .B(_1682_),
    .Y(_1918_));
 sky130_fd_sc_hd__clkinv_4 _3806_ (.A(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__buf_6 _3807_ (.A(_1919_),
    .X(_1132_));
 sky130_fd_sc_hd__a22oi_1 _3808_ (.A1(net382),
    .A2(\stage_gen[4].mux_gen[0].S.IN1_L5 ),
    .B1(net376),
    .B2(\stage_gen[4].mux_gen[0].S.IN1_L3 ),
    .Y(_1920_));
 sky130_fd_sc_hd__nand2_1 _3809_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1384_),
    .Y(_1921_));
 sky130_fd_sc_hd__clkinv_4 _3810_ (.A(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__clkbuf_1 _3811_ (.A(_1922_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _3812_ (.A(net437),
    .B(\stage_gen[5].mux_gen[0].S.IN1_L1 ),
    .Y(_1923_));
 sky130_fd_sc_hd__o21ai_1 _3813_ (.A1(_1917_),
    .A2(_1920_),
    .B1(_1923_),
    .Y(_1208_));
 sky130_fd_sc_hd__clkinv_2 _3814_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .Y(_1924_));
 sky130_fd_sc_hd__and3_1 _3815_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[0].S.IN1_L2 ),
    .X(_1925_));
 sky130_fd_sc_hd__clkbuf_1 _3816_ (.A(_1925_),
    .X(_1210_));
 sky130_fd_sc_hd__nand2b_1 _3817_ (.A_N(_1210_),
    .B(_1923_),
    .Y(_1926_));
 sky130_fd_sc_hd__clkbuf_1 _3818_ (.A(_1926_),
    .X(_1209_));
 sky130_fd_sc_hd__a22oi_2 _3819_ (.A1(net381),
    .A2(\stage_gen[4].mux_gen[1].S.IN1_L5 ),
    .B1(net377),
    .B2(\stage_gen[4].mux_gen[1].S.IN1_L3 ),
    .Y(_1927_));
 sky130_fd_sc_hd__and3_1 _3820_ (.A(_1916_),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[0].S.IN1_L4 ),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _3821_ (.A(_1928_),
    .X(_1212_));
 sky130_fd_sc_hd__o21bai_1 _3822_ (.A1(_1917_),
    .A2(_1927_),
    .B1_N(_1212_),
    .Y(_1211_));
 sky130_fd_sc_hd__a22oi_1 _3823_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[2].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[2].S.IN1_L3 ),
    .Y(_1929_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[1].S.IN1_L1 ),
    .Y(_1930_));
 sky130_fd_sc_hd__o21ai_1 _3825_ (.A1(_1916_),
    .A2(_1929_),
    .B1(_1930_),
    .Y(_1215_));
 sky130_fd_sc_hd__and3_1 _3826_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[1].S.IN1_L2 ),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _3827_ (.A(_1931_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2b_1 _3828_ (.A_N(_1217_),
    .B(_1930_),
    .Y(_1932_));
 sky130_fd_sc_hd__clkbuf_1 _3829_ (.A(_1932_),
    .X(_1216_));
 sky130_fd_sc_hd__a22oi_1 _3830_ (.A1(net385),
    .A2(\stage_gen[4].mux_gen[3].S.IN1_L5 ),
    .B1(net378),
    .B2(\stage_gen[4].mux_gen[3].S.IN1_L3 ),
    .Y(_1933_));
 sky130_fd_sc_hd__and3_1 _3831_ (.A(_1916_),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[1].S.IN1_L4 ),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_1 _3832_ (.A(_1934_),
    .X(_1219_));
 sky130_fd_sc_hd__o21bai_1 _3833_ (.A1(_1917_),
    .A2(_1933_),
    .B1_N(_1219_),
    .Y(_1218_));
 sky130_fd_sc_hd__a22oi_1 _3834_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[4].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[4].S.IN1_L3 ),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[2].S.IN1_L1 ),
    .Y(_1936_));
 sky130_fd_sc_hd__o21ai_1 _3836_ (.A1(_1916_),
    .A2(_1935_),
    .B1(_1936_),
    .Y(_1220_));
 sky130_fd_sc_hd__and3_1 _3837_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[2].S.IN1_L2 ),
    .X(_1937_));
 sky130_fd_sc_hd__clkbuf_1 _3838_ (.A(_1937_),
    .X(_1222_));
 sky130_fd_sc_hd__nand2b_1 _3839_ (.A_N(_1222_),
    .B(_1936_),
    .Y(_1938_));
 sky130_fd_sc_hd__clkbuf_1 _3840_ (.A(_1938_),
    .X(_1221_));
 sky130_fd_sc_hd__a22oi_2 _3841_ (.A1(net386),
    .A2(\stage_gen[4].mux_gen[5].S.IN1_L5 ),
    .B1(net380),
    .B2(\stage_gen[4].mux_gen[5].S.IN1_L3 ),
    .Y(_1939_));
 sky130_fd_sc_hd__and3_1 _3842_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[2].S.IN1_L4 ),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_1 _3843_ (.A(_1940_),
    .X(_1224_));
 sky130_fd_sc_hd__o21bai_1 _3844_ (.A1(_1917_),
    .A2(_1939_),
    .B1_N(_1224_),
    .Y(_1223_));
 sky130_fd_sc_hd__a22oi_1 _3845_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[6].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[6].S.IN1_L3 ),
    .Y(_1941_));
 sky130_fd_sc_hd__nand2_1 _3846_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[3].S.IN1_L1 ),
    .Y(_1942_));
 sky130_fd_sc_hd__o21ai_1 _3847_ (.A1(_1916_),
    .A2(_1941_),
    .B1(_1942_),
    .Y(_1225_));
 sky130_fd_sc_hd__and3_1 _3848_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[3].S.IN1_L2 ),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _3849_ (.A(_1943_),
    .X(_1227_));
 sky130_fd_sc_hd__nand2b_1 _3850_ (.A_N(_1227_),
    .B(_1942_),
    .Y(_1944_));
 sky130_fd_sc_hd__clkbuf_1 _3851_ (.A(_1944_),
    .X(_1226_));
 sky130_fd_sc_hd__a22oi_1 _3852_ (.A1(net385),
    .A2(\stage_gen[4].mux_gen[7].S.IN1_L5 ),
    .B1(net378),
    .B2(\stage_gen[4].mux_gen[7].S.IN1_L3 ),
    .Y(_1945_));
 sky130_fd_sc_hd__and3_1 _3853_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[3].S.IN1_L4 ),
    .X(_1946_));
 sky130_fd_sc_hd__clkbuf_1 _3854_ (.A(_1946_),
    .X(_1229_));
 sky130_fd_sc_hd__o21bai_1 _3855_ (.A1(_1917_),
    .A2(_1945_),
    .B1_N(_1229_),
    .Y(_1228_));
 sky130_fd_sc_hd__a22oi_1 _3856_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[8].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[8].S.IN1_L3 ),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[4].S.IN1_L1 ),
    .Y(_1948_));
 sky130_fd_sc_hd__o21ai_1 _3858_ (.A1(_1916_),
    .A2(_1947_),
    .B1(_1948_),
    .Y(_1230_));
 sky130_fd_sc_hd__and3_1 _3859_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[4].S.IN1_L2 ),
    .X(_1949_));
 sky130_fd_sc_hd__clkbuf_1 _3860_ (.A(_1949_),
    .X(_1232_));
 sky130_fd_sc_hd__nand2b_1 _3861_ (.A_N(_1232_),
    .B(_1948_),
    .Y(_1950_));
 sky130_fd_sc_hd__clkbuf_1 _3862_ (.A(_1950_),
    .X(_1231_));
 sky130_fd_sc_hd__a22oi_1 _3863_ (.A1(net387),
    .A2(\stage_gen[4].mux_gen[9].S.IN1_L5 ),
    .B1(net379),
    .B2(\stage_gen[4].mux_gen[9].S.IN1_L3 ),
    .Y(_1951_));
 sky130_fd_sc_hd__and3_1 _3864_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[4].S.IN1_L4 ),
    .X(_1952_));
 sky130_fd_sc_hd__clkbuf_1 _3865_ (.A(_1952_),
    .X(_1234_));
 sky130_fd_sc_hd__o21bai_1 _3866_ (.A1(_1917_),
    .A2(_1951_),
    .B1_N(_1234_),
    .Y(_1233_));
 sky130_fd_sc_hd__a22oi_1 _3867_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[10].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[10].S.IN1_L3 ),
    .Y(_1953_));
 sky130_fd_sc_hd__nand2_1 _3868_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[5].S.IN1_L1 ),
    .Y(_1954_));
 sky130_fd_sc_hd__o21ai_1 _3869_ (.A1(_1916_),
    .A2(_1953_),
    .B1(_1954_),
    .Y(_1235_));
 sky130_fd_sc_hd__and3_1 _3870_ (.A(_1924_),
    .B(_1892_),
    .C(\stage_gen[5].mux_gen[5].S.IN1_L2 ),
    .X(_1955_));
 sky130_fd_sc_hd__clkbuf_1 _3871_ (.A(_1955_),
    .X(_1237_));
 sky130_fd_sc_hd__nand2b_1 _3872_ (.A_N(_1237_),
    .B(_1954_),
    .Y(_1956_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_1956_),
    .X(_1236_));
 sky130_fd_sc_hd__a22oi_1 _3874_ (.A1(net386),
    .A2(\stage_gen[4].mux_gen[11].S.IN1_L5 ),
    .B1(net379),
    .B2(\stage_gen[4].mux_gen[11].S.IN1_L3 ),
    .Y(_1957_));
 sky130_fd_sc_hd__and3_1 _3875_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1896_),
    .C(\stage_gen[5].mux_gen[5].S.IN1_L4 ),
    .X(_1958_));
 sky130_fd_sc_hd__clkbuf_1 _3876_ (.A(_1958_),
    .X(_1239_));
 sky130_fd_sc_hd__o21bai_1 _3877_ (.A1(_1917_),
    .A2(_1957_),
    .B1_N(_1239_),
    .Y(_1238_));
 sky130_fd_sc_hd__a22oi_1 _3878_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[12].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[12].S.IN1_L3 ),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _3879_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[6].S.IN1_L1 ),
    .Y(_1960_));
 sky130_fd_sc_hd__o21ai_1 _3880_ (.A1(_1916_),
    .A2(_1959_),
    .B1(_1960_),
    .Y(_1240_));
 sky130_fd_sc_hd__buf_6 _3881_ (.A(_1384_),
    .X(_1961_));
 sky130_fd_sc_hd__and3_1 _3882_ (.A(_1924_),
    .B(_1961_),
    .C(\stage_gen[5].mux_gen[6].S.IN1_L2 ),
    .X(_1962_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_1962_),
    .X(_1242_));
 sky130_fd_sc_hd__nand2b_1 _3884_ (.A_N(_1242_),
    .B(_1960_),
    .Y(_1963_));
 sky130_fd_sc_hd__clkbuf_1 _3885_ (.A(_1963_),
    .X(_1241_));
 sky130_fd_sc_hd__a22oi_1 _3886_ (.A1(net382),
    .A2(\stage_gen[4].mux_gen[13].S.IN1_L5 ),
    .B1(net376),
    .B2(\stage_gen[4].mux_gen[13].S.IN1_L3 ),
    .Y(_1964_));
 sky130_fd_sc_hd__buf_4 _3887_ (.A(_1682_),
    .X(_1965_));
 sky130_fd_sc_hd__and3_1 _3888_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1965_),
    .C(\stage_gen[5].mux_gen[6].S.IN1_L4 ),
    .X(_1966_));
 sky130_fd_sc_hd__clkbuf_1 _3889_ (.A(_1966_),
    .X(_1244_));
 sky130_fd_sc_hd__o21bai_1 _3890_ (.A1(_1917_),
    .A2(_1964_),
    .B1_N(_1244_),
    .Y(_1243_));
 sky130_fd_sc_hd__a22oi_1 _3891_ (.A1(_1808_),
    .A2(\stage_gen[4].mux_gen[14].S.IN1_L5 ),
    .B1(_1919_),
    .B2(\stage_gen[4].mux_gen[14].S.IN1_L3 ),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _3892_ (.A(_1922_),
    .B(\stage_gen[5].mux_gen[7].S.IN1_L1 ),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_1 _3893_ (.A1(_1916_),
    .A2(_1967_),
    .B1(_1968_),
    .Y(_1245_));
 sky130_fd_sc_hd__and3_1 _3894_ (.A(_1924_),
    .B(_1961_),
    .C(\stage_gen[5].mux_gen[7].S.IN1_L2 ),
    .X(_1969_));
 sky130_fd_sc_hd__clkbuf_1 _3895_ (.A(_1969_),
    .X(_1247_));
 sky130_fd_sc_hd__nand2b_1 _3896_ (.A_N(_1247_),
    .B(_1968_),
    .Y(_1970_));
 sky130_fd_sc_hd__clkbuf_1 _3897_ (.A(_1970_),
    .X(_1246_));
 sky130_fd_sc_hd__a22oi_1 _3898_ (.A1(net381),
    .A2(\stage_gen[4].mux_gen[15].S.IN1_L5 ),
    .B1(net376),
    .B2(\stage_gen[4].mux_gen[15].S.IN1_L3 ),
    .Y(_1971_));
 sky130_fd_sc_hd__and3_1 _3899_ (.A(\stage_gen[5].genblk1.clks.clk_o ),
    .B(_1965_),
    .C(\stage_gen[5].mux_gen[7].S.IN1_L4 ),
    .X(_1972_));
 sky130_fd_sc_hd__clkbuf_1 _3900_ (.A(_1972_),
    .X(_1249_));
 sky130_fd_sc_hd__o21bai_1 _3901_ (.A1(_1917_),
    .A2(_1971_),
    .B1_N(_1249_),
    .Y(_1248_));
 sky130_fd_sc_hd__buf_2 _3902_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .X(_1973_));
 sky130_fd_sc_hd__nand2_1 _3903_ (.A(_1924_),
    .B(_1801_),
    .Y(_1974_));
 sky130_fd_sc_hd__clkinv_4 _3904_ (.A(_1974_),
    .Y(_1214_));
 sky130_fd_sc_hd__a22oi_1 _3905_ (.A1(net437),
    .A2(\stage_gen[5].mux_gen[0].S.IN1_L5 ),
    .B1(net435),
    .B2(\stage_gen[5].mux_gen[0].S.IN1_L3 ),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .B(_1801_),
    .Y(_1976_));
 sky130_fd_sc_hd__clkinv_4 _3907_ (.A(_1976_),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(net433),
    .B(\stage_gen[6].mux_gen[0].S.IN1_L1 ),
    .Y(_1977_));
 sky130_fd_sc_hd__o21ai_1 _3909_ (.A1(_1973_),
    .A2(_1975_),
    .B1(_1977_),
    .Y(_1250_));
 sky130_fd_sc_hd__inv_2 _3910_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .Y(_1978_));
 sky130_fd_sc_hd__and3_1 _3911_ (.A(_1978_),
    .B(_1961_),
    .C(\stage_gen[6].mux_gen[0].S.IN1_L2 ),
    .X(_1979_));
 sky130_fd_sc_hd__clkbuf_1 _3912_ (.A(_1979_),
    .X(_1252_));
 sky130_fd_sc_hd__or2b_1 _3913_ (.A(_1252_),
    .B_N(_1977_),
    .X(_1980_));
 sky130_fd_sc_hd__clkbuf_1 _3914_ (.A(_1980_),
    .X(_1251_));
 sky130_fd_sc_hd__a22oi_1 _3915_ (.A1(net439),
    .A2(\stage_gen[5].mux_gen[1].S.IN1_L5 ),
    .B1(net435),
    .B2(\stage_gen[5].mux_gen[1].S.IN1_L3 ),
    .Y(_1981_));
 sky130_fd_sc_hd__and3_1 _3916_ (.A(_1973_),
    .B(_1965_),
    .C(\stage_gen[6].mux_gen[0].S.IN1_L4 ),
    .X(_1982_));
 sky130_fd_sc_hd__clkbuf_1 _3917_ (.A(_1982_),
    .X(_1254_));
 sky130_fd_sc_hd__o21bai_1 _3918_ (.A1(_1973_),
    .A2(_1981_),
    .B1_N(_1254_),
    .Y(_1253_));
 sky130_fd_sc_hd__a22oi_1 _3919_ (.A1(net439),
    .A2(\stage_gen[5].mux_gen[2].S.IN1_L5 ),
    .B1(net434),
    .B2(\stage_gen[5].mux_gen[2].S.IN1_L3 ),
    .Y(_1983_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(net433),
    .B(\stage_gen[6].mux_gen[1].S.IN1_L1 ),
    .Y(_1984_));
 sky130_fd_sc_hd__o21ai_1 _3921_ (.A1(_1973_),
    .A2(_1983_),
    .B1(_1984_),
    .Y(_1257_));
 sky130_fd_sc_hd__and3_1 _3922_ (.A(_1978_),
    .B(_1961_),
    .C(\stage_gen[6].mux_gen[1].S.IN1_L2 ),
    .X(_1985_));
 sky130_fd_sc_hd__clkbuf_1 _3923_ (.A(_1985_),
    .X(_1259_));
 sky130_fd_sc_hd__or2b_1 _3924_ (.A(_1259_),
    .B_N(_1984_),
    .X(_1986_));
 sky130_fd_sc_hd__clkbuf_1 _3925_ (.A(_1986_),
    .X(_1258_));
 sky130_fd_sc_hd__a22oi_1 _3926_ (.A1(net439),
    .A2(\stage_gen[5].mux_gen[3].S.IN1_L5 ),
    .B1(net434),
    .B2(\stage_gen[5].mux_gen[3].S.IN1_L3 ),
    .Y(_1987_));
 sky130_fd_sc_hd__and3_1 _3927_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .B(_1965_),
    .C(\stage_gen[6].mux_gen[1].S.IN1_L4 ),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_1 _3928_ (.A(_1988_),
    .X(_1261_));
 sky130_fd_sc_hd__o21bai_1 _3929_ (.A1(_1973_),
    .A2(_1987_),
    .B1_N(_1261_),
    .Y(_1260_));
 sky130_fd_sc_hd__a22oi_1 _3930_ (.A1(net439),
    .A2(\stage_gen[5].mux_gen[4].S.IN1_L5 ),
    .B1(net434),
    .B2(\stage_gen[5].mux_gen[4].S.IN1_L3 ),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(net433),
    .B(\stage_gen[6].mux_gen[2].S.IN1_L1 ),
    .Y(_1990_));
 sky130_fd_sc_hd__o21ai_1 _3932_ (.A1(_1973_),
    .A2(_1989_),
    .B1(_1990_),
    .Y(_1262_));
 sky130_fd_sc_hd__and3_1 _3933_ (.A(_1978_),
    .B(_1961_),
    .C(\stage_gen[6].mux_gen[2].S.IN1_L2 ),
    .X(_1991_));
 sky130_fd_sc_hd__clkbuf_1 _3934_ (.A(_1991_),
    .X(_1264_));
 sky130_fd_sc_hd__or2b_1 _3935_ (.A(_1264_),
    .B_N(_1990_),
    .X(_1992_));
 sky130_fd_sc_hd__clkbuf_1 _3936_ (.A(_1992_),
    .X(_1263_));
 sky130_fd_sc_hd__a22oi_1 _3937_ (.A1(net439),
    .A2(\stage_gen[5].mux_gen[5].S.IN1_L5 ),
    .B1(net434),
    .B2(\stage_gen[5].mux_gen[5].S.IN1_L3 ),
    .Y(_1993_));
 sky130_fd_sc_hd__and3_1 _3938_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .B(_1965_),
    .C(\stage_gen[6].mux_gen[2].S.IN1_L4 ),
    .X(_1994_));
 sky130_fd_sc_hd__clkbuf_1 _3939_ (.A(_1994_),
    .X(_1266_));
 sky130_fd_sc_hd__o21bai_1 _3940_ (.A1(_1973_),
    .A2(_1993_),
    .B1_N(_1266_),
    .Y(_1265_));
 sky130_fd_sc_hd__a22oi_1 _3941_ (.A1(net437),
    .A2(\stage_gen[5].mux_gen[6].S.IN1_L5 ),
    .B1(net435),
    .B2(\stage_gen[5].mux_gen[6].S.IN1_L3 ),
    .Y(_1995_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(net432),
    .B(\stage_gen[6].mux_gen[3].S.IN1_L1 ),
    .Y(_1996_));
 sky130_fd_sc_hd__o21ai_1 _3943_ (.A1(_1973_),
    .A2(_1995_),
    .B1(_1996_),
    .Y(_1267_));
 sky130_fd_sc_hd__and3_1 _3944_ (.A(_1978_),
    .B(_1961_),
    .C(\stage_gen[6].mux_gen[3].S.IN1_L2 ),
    .X(_1997_));
 sky130_fd_sc_hd__clkbuf_1 _3945_ (.A(_1997_),
    .X(_1269_));
 sky130_fd_sc_hd__or2b_1 _3946_ (.A(_1269_),
    .B_N(_1996_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_1 _3947_ (.A(_1998_),
    .X(_1268_));
 sky130_fd_sc_hd__a22oi_1 _3948_ (.A1(net437),
    .A2(\stage_gen[5].mux_gen[7].S.IN1_L5 ),
    .B1(net435),
    .B2(\stage_gen[5].mux_gen[7].S.IN1_L3 ),
    .Y(_1999_));
 sky130_fd_sc_hd__and3_1 _3949_ (.A(\stage_gen[6].genblk1.clks.clk_o ),
    .B(_1965_),
    .C(\stage_gen[6].mux_gen[3].S.IN1_L4 ),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _3950_ (.A(_2000_),
    .X(_1271_));
 sky130_fd_sc_hd__o21bai_1 _3951_ (.A1(_1973_),
    .A2(_1999_),
    .B1_N(_1271_),
    .Y(_1270_));
 sky130_fd_sc_hd__buf_2 _3952_ (.A(\stage_gen[7].genblk1.clks.clk_o ),
    .X(_2001_));
 sky130_fd_sc_hd__nand2_1 _3953_ (.A(_1978_),
    .B(_1801_),
    .Y(_2002_));
 sky130_fd_sc_hd__inv_2 _3954_ (.A(_2002_),
    .Y(_1256_));
 sky130_fd_sc_hd__a22oi_1 _3955_ (.A1(net433),
    .A2(\stage_gen[6].mux_gen[0].S.IN1_L5 ),
    .B1(_1256_),
    .B2(\stage_gen[6].mux_gen[0].S.IN1_L3 ),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _3956_ (.A(_2001_),
    .B(_1377_),
    .Y(_2004_));
 sky130_fd_sc_hd__clkinv_2 _3957_ (.A(_2004_),
    .Y(_1277_));
 sky130_fd_sc_hd__nand2_1 _3958_ (.A(_1277_),
    .B(\stage_gen[7].mux_gen[0].S.IN1_L1 ),
    .Y(_2005_));
 sky130_fd_sc_hd__o21ai_1 _3959_ (.A1(_2001_),
    .A2(_2003_),
    .B1(_2005_),
    .Y(_1272_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(_2001_),
    .Y(_2006_));
 sky130_fd_sc_hd__and3_1 _3961_ (.A(_2006_),
    .B(_1961_),
    .C(\stage_gen[7].mux_gen[0].S.IN1_L2 ),
    .X(_2007_));
 sky130_fd_sc_hd__clkbuf_1 _3962_ (.A(_2007_),
    .X(_1274_));
 sky130_fd_sc_hd__nand2b_1 _3963_ (.A_N(_1274_),
    .B(_2005_),
    .Y(_2008_));
 sky130_fd_sc_hd__clkbuf_1 _3964_ (.A(_2008_),
    .X(_1273_));
 sky130_fd_sc_hd__a22oi_1 _3965_ (.A1(net433),
    .A2(\stage_gen[6].mux_gen[1].S.IN1_L5 ),
    .B1(net431),
    .B2(\stage_gen[6].mux_gen[1].S.IN1_L3 ),
    .Y(_2009_));
 sky130_fd_sc_hd__and3_1 _3966_ (.A(_2001_),
    .B(_1965_),
    .C(\stage_gen[7].mux_gen[0].S.IN1_L4 ),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _3967_ (.A(_2010_),
    .X(_1276_));
 sky130_fd_sc_hd__o21bai_1 _3968_ (.A1(_2001_),
    .A2(_2009_),
    .B1_N(_1276_),
    .Y(_1275_));
 sky130_fd_sc_hd__a22oi_1 _3969_ (.A1(net432),
    .A2(\stage_gen[6].mux_gen[2].S.IN1_L5 ),
    .B1(net431),
    .B2(\stage_gen[6].mux_gen[2].S.IN1_L3 ),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_1277_),
    .B(\stage_gen[7].mux_gen[1].S.IN1_L1 ),
    .Y(_2012_));
 sky130_fd_sc_hd__o21ai_1 _3971_ (.A1(_2001_),
    .A2(_2011_),
    .B1(_2012_),
    .Y(_1279_));
 sky130_fd_sc_hd__and3_1 _3972_ (.A(_2006_),
    .B(_1961_),
    .C(\stage_gen[7].mux_gen[1].S.IN1_L2 ),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _3973_ (.A(_2013_),
    .X(_1281_));
 sky130_fd_sc_hd__nand2b_1 _3974_ (.A_N(_1281_),
    .B(_2012_),
    .Y(_2014_));
 sky130_fd_sc_hd__clkbuf_1 _3975_ (.A(_2014_),
    .X(_1280_));
 sky130_fd_sc_hd__a22oi_1 _3976_ (.A1(net432),
    .A2(\stage_gen[6].mux_gen[3].S.IN1_L5 ),
    .B1(net431),
    .B2(\stage_gen[6].mux_gen[3].S.IN1_L3 ),
    .Y(_2015_));
 sky130_fd_sc_hd__and3_1 _3977_ (.A(_2001_),
    .B(_1965_),
    .C(\stage_gen[7].mux_gen[1].S.IN1_L4 ),
    .X(_2016_));
 sky130_fd_sc_hd__clkbuf_1 _3978_ (.A(_2016_),
    .X(_1283_));
 sky130_fd_sc_hd__o21bai_1 _3979_ (.A1(_2001_),
    .A2(_2015_),
    .B1_N(_1283_),
    .Y(_1282_));
 sky130_fd_sc_hd__buf_4 _3980_ (.A(clknet_3_2__leaf_CLK),
    .X(_2017_));
 sky130_fd_sc_hd__buf_2 _3981_ (.A(clknet_1_0__leaf__2017_),
    .X(_2018_));
 sky130_fd_sc_hd__buf_4 _3982_ (.A(_1390_),
    .X(_2019_));
 sky130_fd_sc_hd__nand2_1 _3983_ (.A(_2006_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__inv_2 _3984_ (.A(_2020_),
    .Y(_1278_));
 sky130_fd_sc_hd__a22oi_1 _3985_ (.A1(_1277_),
    .A2(\stage_gen[7].mux_gen[0].S.IN1_L5 ),
    .B1(_1278_),
    .B2(\stage_gen[7].mux_gen[0].S.IN1_L3 ),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_4 _3986_ (.A(clknet_1_1__leaf__2017_),
    .B(_1361_),
    .Y(_2022_));
 sky130_fd_sc_hd__inv_4 _3987__13 (.A(clknet_1_0__leaf__2022_),
    .Y(net453));
 sky130_fd_sc_hd__inv_4 _3987__14 (.A(clknet_1_1__leaf__2022_),
    .Y(net454));
 sky130_fd_sc_hd__inv_4 _3987__15 (.A(clknet_1_1__leaf__2022_),
    .Y(net455));
 sky130_fd_sc_hd__inv_4 _3987__16 (.A(clknet_1_0__leaf__2022_),
    .Y(net456));
 sky130_fd_sc_hd__inv_4 _3987__17 (.A(clknet_1_1__leaf__2022_),
    .Y(net457));
 sky130_fd_sc_hd__inv_4 _3987__18 (.A(clknet_1_0__leaf__2022_),
    .Y(net458));
 sky130_fd_sc_hd__inv_4 _3987__19 (.A(clknet_1_0__leaf__2022_),
    .Y(net459));
 sky130_fd_sc_hd__inv_4 _3987__20 (.A(clknet_1_0__leaf__2022_),
    .Y(net460));
 sky130_fd_sc_hd__inv_4 _3987__21 (.A(clknet_1_0__leaf__2022_),
    .Y(net461));
 sky130_fd_sc_hd__inv_4 _3987__22 (.A(clknet_1_1__leaf__2022_),
    .Y(net462));
 sky130_fd_sc_hd__nand2_2 _3988_ (.A(net462),
    .B(\stage_gen[8].mux_gen[0].S.IN1_L1 ),
    .Y(_2023_));
 sky130_fd_sc_hd__o21ai_2 _3989_ (.A1(clknet_1_1__leaf__2018_),
    .A2(_2021_),
    .B1(clknet_1_1__leaf__2023_),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _3990__1 (.A(clknet_3_5__leaf_CLK),
    .Y(net441));
 sky130_fd_sc_hd__and3_4 _3991_ (.A(net444),
    .B(_1961_),
    .C(\stage_gen[8].mux_gen[0].S.IN1_L2 ),
    .X(_2025_));
 sky130_fd_sc_hd__buf_6 _3992_ (.A(_2025_),
    .X(_1286_));
 sky130_fd_sc_hd__nand2b_4 _3993_ (.A_N(clknet_1_1__leaf__1286_),
    .B(clknet_1_0__leaf__2023_),
    .Y(_2026_));
 sky130_fd_sc_hd__buf_6 _3994_ (.A(_2026_),
    .X(_1285_));
 sky130_fd_sc_hd__inv_2 _3995_ (.A(\stage_gen[8].mux_gen[0].S.IN1_L4 ),
    .Y(_2027_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(\stage_gen[7].mux_gen[1].S.IN1_L3 ),
    .A1(\stage_gen[7].mux_gen[1].S.IN1_L5 ),
    .S(_2001_),
    .X(_2028_));
 sky130_fd_sc_hd__buf_4 _3997_ (.A(_2019_),
    .X(_2029_));
 sky130_fd_sc_hd__nand3_2 _3998_ (.A(_2028_),
    .B(net443),
    .C(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__o21ai_2 _3999_ (.A1(_2027_),
    .A2(clknet_1_1__leaf__2022_),
    .B1(_2030_),
    .Y(_1287_));
 sky130_fd_sc_hd__mux2_2 _4000_ (.A0(\stage_gen[8].mux_gen[0].S.IN1_L3 ),
    .A1(\stage_gen[8].mux_gen[0].S.IN1_L5 ),
    .S(clknet_1_1__leaf__2017_),
    .X(_2031_));
 sky130_fd_sc_hd__buf_1 _4001_ (.A(_2031_),
    .X(net258));
 sky130_fd_sc_hd__buf_4 _4002_ (.A(_1373_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _4003_ (.A(_2032_),
    .X(_0006_));
 sky130_fd_sc_hd__clkbuf_4 _4004_ (.A(_1368_),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_2 _4005_ (.A(_2033_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_4 _4006_ (.A(\stage_gen[1].genblk1.clks.clk_o ),
    .X(_2034_));
 sky130_fd_sc_hd__and3_1 _4007_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[0].S.IN1_L4 ),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _4008_ (.A(_2035_),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _4009_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[1].S.IN1_L4 ),
    .X(_2036_));
 sky130_fd_sc_hd__clkbuf_1 _4010_ (.A(_2036_),
    .X(_0201_));
 sky130_fd_sc_hd__and3_1 _4011_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[2].S.IN1_L4 ),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _4012_ (.A(_2037_),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[3].S.IN1_L4 ),
    .X(_2038_));
 sky130_fd_sc_hd__clkbuf_1 _4014_ (.A(_2038_),
    .X(_0311_));
 sky130_fd_sc_hd__and3_1 _4015_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[4].S.IN1_L4 ),
    .X(_2039_));
 sky130_fd_sc_hd__clkbuf_1 _4016_ (.A(_2039_),
    .X(_0366_));
 sky130_fd_sc_hd__and3_1 _4017_ (.A(_2034_),
    .B(_2019_),
    .C(\stage_gen[1].mux_gen[5].S.IN1_L4 ),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_1 _4018_ (.A(_2040_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_6 _4019_ (.A(_1360_),
    .X(_2041_));
 sky130_fd_sc_hd__buf_2 _4020_ (.A(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__and3_1 _4021_ (.A(_2034_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[6].S.IN1_L4 ),
    .X(_2043_));
 sky130_fd_sc_hd__clkbuf_1 _4022_ (.A(_2043_),
    .X(_0476_));
 sky130_fd_sc_hd__and3_1 _4023_ (.A(_2034_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[7].S.IN1_L4 ),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _4024_ (.A(_2044_),
    .X(_0531_));
 sky130_fd_sc_hd__and3_1 _4025_ (.A(_2034_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[8].S.IN1_L4 ),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _4026_ (.A(_2045_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_4 _4027_ (.A(\stage_gen[1].genblk1.clks.clk_o ),
    .X(_2046_));
 sky130_fd_sc_hd__buf_2 _4028_ (.A(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__and3_1 _4029_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[9].S.IN1_L4 ),
    .X(_2048_));
 sky130_fd_sc_hd__clkbuf_1 _4030_ (.A(_2048_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _4031_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[10].S.IN1_L4 ),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _4032_ (.A(_2049_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _4033_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[11].S.IN1_L4 ),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _4034_ (.A(_2050_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _4035_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[12].S.IN1_L4 ),
    .X(_2051_));
 sky130_fd_sc_hd__clkbuf_1 _4036_ (.A(_2051_),
    .X(_0161_));
 sky130_fd_sc_hd__and3_1 _4037_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[13].S.IN1_L4 ),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _4038_ (.A(_2052_),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _4039_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[14].S.IN1_L4 ),
    .X(_2053_));
 sky130_fd_sc_hd__clkbuf_1 _4040_ (.A(_2053_),
    .X(_0171_));
 sky130_fd_sc_hd__and3_1 _4041_ (.A(_2047_),
    .B(_2042_),
    .C(\stage_gen[1].mux_gen[15].S.IN1_L4 ),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _4042_ (.A(_2054_),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_4 _4043_ (.A(_2041_),
    .X(_2055_));
 sky130_fd_sc_hd__and3_1 _4044_ (.A(_2047_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[16].S.IN1_L4 ),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _4045_ (.A(_2056_),
    .X(_0181_));
 sky130_fd_sc_hd__and3_1 _4046_ (.A(_2047_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[17].S.IN1_L4 ),
    .X(_2057_));
 sky130_fd_sc_hd__clkbuf_1 _4047_ (.A(_2057_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _4048_ (.A(_2047_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[18].S.IN1_L4 ),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _4049_ (.A(_2058_),
    .X(_0191_));
 sky130_fd_sc_hd__buf_4 _4050_ (.A(\stage_gen[1].genblk1.clks.clk_o ),
    .X(_2059_));
 sky130_fd_sc_hd__buf_2 _4051_ (.A(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__and3_1 _4052_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[19].S.IN1_L4 ),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_1 _4053_ (.A(_2061_),
    .X(_0196_));
 sky130_fd_sc_hd__and3_1 _4054_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[20].S.IN1_L4 ),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _4055_ (.A(_2062_),
    .X(_0206_));
 sky130_fd_sc_hd__and3_1 _4056_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[21].S.IN1_L4 ),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _4057_ (.A(_2063_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_1 _4058_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[22].S.IN1_L4 ),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _4059_ (.A(_2064_),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _4060_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[23].S.IN1_L4 ),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _4061_ (.A(_2065_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _4062_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[24].S.IN1_L4 ),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _4063_ (.A(_2066_),
    .X(_0226_));
 sky130_fd_sc_hd__and3_1 _4064_ (.A(_2060_),
    .B(_2055_),
    .C(\stage_gen[1].mux_gen[25].S.IN1_L4 ),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_1 _4065_ (.A(_2067_),
    .X(_0231_));
 sky130_fd_sc_hd__buf_2 _4066_ (.A(_2041_),
    .X(_2068_));
 sky130_fd_sc_hd__and3_1 _4067_ (.A(_2060_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[26].S.IN1_L4 ),
    .X(_2069_));
 sky130_fd_sc_hd__clkbuf_1 _4068_ (.A(_2069_),
    .X(_0236_));
 sky130_fd_sc_hd__and3_1 _4069_ (.A(_2060_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[27].S.IN1_L4 ),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _4070_ (.A(_2070_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _4071_ (.A(_2060_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[28].S.IN1_L4 ),
    .X(_2071_));
 sky130_fd_sc_hd__clkbuf_1 _4072_ (.A(_2071_),
    .X(_0246_));
 sky130_fd_sc_hd__buf_2 _4073_ (.A(_2059_),
    .X(_2072_));
 sky130_fd_sc_hd__and3_1 _4074_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[29].S.IN1_L4 ),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_1 _4075_ (.A(_2073_),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _4076_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[30].S.IN1_L4 ),
    .X(_2074_));
 sky130_fd_sc_hd__clkbuf_1 _4077_ (.A(_2074_),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _4078_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[31].S.IN1_L4 ),
    .X(_2075_));
 sky130_fd_sc_hd__clkbuf_1 _4079_ (.A(_2075_),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _4080_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[32].S.IN1_L4 ),
    .X(_2076_));
 sky130_fd_sc_hd__clkbuf_1 _4081_ (.A(_2076_),
    .X(_0271_));
 sky130_fd_sc_hd__and3_1 _4082_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[33].S.IN1_L4 ),
    .X(_2077_));
 sky130_fd_sc_hd__clkbuf_1 _4083_ (.A(_2077_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _4084_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[34].S.IN1_L4 ),
    .X(_2078_));
 sky130_fd_sc_hd__clkbuf_1 _4085_ (.A(_2078_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _4086_ (.A(_2072_),
    .B(_2068_),
    .C(\stage_gen[1].mux_gen[35].S.IN1_L4 ),
    .X(_2079_));
 sky130_fd_sc_hd__clkbuf_1 _4087_ (.A(_2079_),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _4088_ (.A(_2041_),
    .X(_2080_));
 sky130_fd_sc_hd__and3_1 _4089_ (.A(_2072_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[36].S.IN1_L4 ),
    .X(_2081_));
 sky130_fd_sc_hd__clkbuf_1 _4090_ (.A(_2081_),
    .X(_0291_));
 sky130_fd_sc_hd__and3_1 _4091_ (.A(_2072_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[37].S.IN1_L4 ),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _4092_ (.A(_2082_),
    .X(_0296_));
 sky130_fd_sc_hd__and3_1 _4093_ (.A(_2072_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[38].S.IN1_L4 ),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _4094_ (.A(_2083_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_2 _4095_ (.A(_2059_),
    .X(_2084_));
 sky130_fd_sc_hd__and3_1 _4096_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[39].S.IN1_L4 ),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_1 _4097_ (.A(_2085_),
    .X(_0306_));
 sky130_fd_sc_hd__and3_1 _4098_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[40].S.IN1_L4 ),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _4099_ (.A(_2086_),
    .X(_0316_));
 sky130_fd_sc_hd__and3_1 _4100_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[41].S.IN1_L4 ),
    .X(_2087_));
 sky130_fd_sc_hd__clkbuf_1 _4101_ (.A(_2087_),
    .X(_0321_));
 sky130_fd_sc_hd__and3_1 _4102_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[42].S.IN1_L4 ),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_1 _4103_ (.A(_2088_),
    .X(_0326_));
 sky130_fd_sc_hd__and3_1 _4104_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[43].S.IN1_L4 ),
    .X(_2089_));
 sky130_fd_sc_hd__clkbuf_1 _4105_ (.A(_2089_),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _4106_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[44].S.IN1_L4 ),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_1 _4107_ (.A(_2090_),
    .X(_0336_));
 sky130_fd_sc_hd__and3_1 _4108_ (.A(_2084_),
    .B(_2080_),
    .C(\stage_gen[1].mux_gen[45].S.IN1_L4 ),
    .X(_2091_));
 sky130_fd_sc_hd__clkbuf_1 _4109_ (.A(_2091_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_2 _4110_ (.A(_2041_),
    .X(_2092_));
 sky130_fd_sc_hd__and3_1 _4111_ (.A(_2084_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[46].S.IN1_L4 ),
    .X(_2093_));
 sky130_fd_sc_hd__clkbuf_1 _4112_ (.A(_2093_),
    .X(_0346_));
 sky130_fd_sc_hd__and3_1 _4113_ (.A(_2084_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[47].S.IN1_L4 ),
    .X(_2094_));
 sky130_fd_sc_hd__clkbuf_1 _4114_ (.A(_2094_),
    .X(_0351_));
 sky130_fd_sc_hd__and3_1 _4115_ (.A(_2084_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[48].S.IN1_L4 ),
    .X(_2095_));
 sky130_fd_sc_hd__clkbuf_1 _4116_ (.A(_2095_),
    .X(_0356_));
 sky130_fd_sc_hd__buf_2 _4117_ (.A(_2059_),
    .X(_2096_));
 sky130_fd_sc_hd__and3_1 _4118_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[49].S.IN1_L4 ),
    .X(_2097_));
 sky130_fd_sc_hd__clkbuf_1 _4119_ (.A(_2097_),
    .X(_0361_));
 sky130_fd_sc_hd__and3_1 _4120_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[50].S.IN1_L4 ),
    .X(_2098_));
 sky130_fd_sc_hd__clkbuf_1 _4121_ (.A(_2098_),
    .X(_0371_));
 sky130_fd_sc_hd__and3_1 _4122_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[51].S.IN1_L4 ),
    .X(_2099_));
 sky130_fd_sc_hd__clkbuf_1 _4123_ (.A(_2099_),
    .X(_0376_));
 sky130_fd_sc_hd__and3_1 _4124_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[52].S.IN1_L4 ),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_1 _4125_ (.A(_2100_),
    .X(_0381_));
 sky130_fd_sc_hd__and3_1 _4126_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[53].S.IN1_L4 ),
    .X(_2101_));
 sky130_fd_sc_hd__clkbuf_1 _4127_ (.A(_2101_),
    .X(_0386_));
 sky130_fd_sc_hd__and3_1 _4128_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[54].S.IN1_L4 ),
    .X(_2102_));
 sky130_fd_sc_hd__clkbuf_1 _4129_ (.A(_2102_),
    .X(_0391_));
 sky130_fd_sc_hd__and3_1 _4130_ (.A(_2096_),
    .B(_2092_),
    .C(\stage_gen[1].mux_gen[55].S.IN1_L4 ),
    .X(_2103_));
 sky130_fd_sc_hd__clkbuf_1 _4131_ (.A(_2103_),
    .X(_0396_));
 sky130_fd_sc_hd__buf_2 _4132_ (.A(_2041_),
    .X(_2104_));
 sky130_fd_sc_hd__and3_1 _4133_ (.A(_2096_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[56].S.IN1_L4 ),
    .X(_2105_));
 sky130_fd_sc_hd__clkbuf_1 _4134_ (.A(_2105_),
    .X(_0401_));
 sky130_fd_sc_hd__and3_1 _4135_ (.A(_2096_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[57].S.IN1_L4 ),
    .X(_2106_));
 sky130_fd_sc_hd__clkbuf_1 _4136_ (.A(_2106_),
    .X(_0406_));
 sky130_fd_sc_hd__and3_1 _4137_ (.A(_2096_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[58].S.IN1_L4 ),
    .X(_2107_));
 sky130_fd_sc_hd__clkbuf_1 _4138_ (.A(_2107_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_2 _4139_ (.A(_2059_),
    .X(_2108_));
 sky130_fd_sc_hd__and3_1 _4140_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[59].S.IN1_L4 ),
    .X(_2109_));
 sky130_fd_sc_hd__clkbuf_1 _4141_ (.A(_2109_),
    .X(_0416_));
 sky130_fd_sc_hd__and3_1 _4142_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[60].S.IN1_L4 ),
    .X(_2110_));
 sky130_fd_sc_hd__clkbuf_1 _4143_ (.A(_2110_),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _4144_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[61].S.IN1_L4 ),
    .X(_2111_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_2111_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _4146_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[62].S.IN1_L4 ),
    .X(_2112_));
 sky130_fd_sc_hd__clkbuf_1 _4147_ (.A(_2112_),
    .X(_0436_));
 sky130_fd_sc_hd__and3_1 _4148_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[63].S.IN1_L4 ),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_2113_),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _4150_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[64].S.IN1_L4 ),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_1 _4151_ (.A(_2114_),
    .X(_0446_));
 sky130_fd_sc_hd__and3_1 _4152_ (.A(_2108_),
    .B(_2104_),
    .C(\stage_gen[1].mux_gen[65].S.IN1_L4 ),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_2115_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _4154_ (.A(_2041_),
    .X(_2116_));
 sky130_fd_sc_hd__and3_1 _4155_ (.A(_2108_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[66].S.IN1_L4 ),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _4156_ (.A(_2117_),
    .X(_0456_));
 sky130_fd_sc_hd__and3_1 _4157_ (.A(_2108_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[67].S.IN1_L4 ),
    .X(_2118_));
 sky130_fd_sc_hd__clkbuf_1 _4158_ (.A(_2118_),
    .X(_0461_));
 sky130_fd_sc_hd__and3_1 _4159_ (.A(_2108_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[68].S.IN1_L4 ),
    .X(_2119_));
 sky130_fd_sc_hd__clkbuf_1 _4160_ (.A(_2119_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _4161_ (.A(_2059_),
    .X(_2120_));
 sky130_fd_sc_hd__and3_1 _4162_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[69].S.IN1_L4 ),
    .X(_2121_));
 sky130_fd_sc_hd__clkbuf_1 _4163_ (.A(_2121_),
    .X(_0471_));
 sky130_fd_sc_hd__and3_1 _4164_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[70].S.IN1_L4 ),
    .X(_2122_));
 sky130_fd_sc_hd__clkbuf_1 _4165_ (.A(_2122_),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _4166_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[71].S.IN1_L4 ),
    .X(_2123_));
 sky130_fd_sc_hd__clkbuf_1 _4167_ (.A(_2123_),
    .X(_0486_));
 sky130_fd_sc_hd__and3_1 _4168_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[72].S.IN1_L4 ),
    .X(_2124_));
 sky130_fd_sc_hd__clkbuf_1 _4169_ (.A(_2124_),
    .X(_0491_));
 sky130_fd_sc_hd__and3_1 _4170_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[73].S.IN1_L4 ),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_1 _4171_ (.A(_2125_),
    .X(_0496_));
 sky130_fd_sc_hd__and3_1 _4172_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[74].S.IN1_L4 ),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_1 _4173_ (.A(_2126_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _4174_ (.A(_2120_),
    .B(_2116_),
    .C(\stage_gen[1].mux_gen[75].S.IN1_L4 ),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_1 _4175_ (.A(_2127_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_4 _4176_ (.A(_2041_),
    .X(_2128_));
 sky130_fd_sc_hd__and3_1 _4177_ (.A(_2120_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[76].S.IN1_L4 ),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _4178_ (.A(_2129_),
    .X(_0511_));
 sky130_fd_sc_hd__and3_1 _4179_ (.A(_2120_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[77].S.IN1_L4 ),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _4180_ (.A(_2130_),
    .X(_0516_));
 sky130_fd_sc_hd__and3_1 _4181_ (.A(_2120_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[78].S.IN1_L4 ),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _4182_ (.A(_2131_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _4183_ (.A(_2059_),
    .X(_2132_));
 sky130_fd_sc_hd__and3_1 _4184_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[79].S.IN1_L4 ),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _4185_ (.A(_2133_),
    .X(_0526_));
 sky130_fd_sc_hd__and3_1 _4186_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[80].S.IN1_L4 ),
    .X(_2134_));
 sky130_fd_sc_hd__clkbuf_1 _4187_ (.A(_2134_),
    .X(_0536_));
 sky130_fd_sc_hd__and3_1 _4188_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[81].S.IN1_L4 ),
    .X(_2135_));
 sky130_fd_sc_hd__clkbuf_1 _4189_ (.A(_2135_),
    .X(_0541_));
 sky130_fd_sc_hd__and3_1 _4190_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[82].S.IN1_L4 ),
    .X(_2136_));
 sky130_fd_sc_hd__clkbuf_1 _4191_ (.A(_2136_),
    .X(_0546_));
 sky130_fd_sc_hd__and3_1 _4192_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[83].S.IN1_L4 ),
    .X(_2137_));
 sky130_fd_sc_hd__clkbuf_1 _4193_ (.A(_2137_),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _4194_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[84].S.IN1_L4 ),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_1 _4195_ (.A(_2138_),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _4196_ (.A(_2132_),
    .B(_2128_),
    .C(\stage_gen[1].mux_gen[85].S.IN1_L4 ),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_1 _4197_ (.A(_2139_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_4 _4198_ (.A(_2041_),
    .X(_2140_));
 sky130_fd_sc_hd__and3_1 _4199_ (.A(_2132_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[86].S.IN1_L4 ),
    .X(_2141_));
 sky130_fd_sc_hd__clkbuf_1 _4200_ (.A(_2141_),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _4201_ (.A(_2132_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[87].S.IN1_L4 ),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _4202_ (.A(_2142_),
    .X(_0571_));
 sky130_fd_sc_hd__and3_1 _4203_ (.A(_2132_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[88].S.IN1_L4 ),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_1 _4204_ (.A(_2143_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_4 _4205_ (.A(_2059_),
    .X(_2144_));
 sky130_fd_sc_hd__and3_1 _4206_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[89].S.IN1_L4 ),
    .X(_2145_));
 sky130_fd_sc_hd__clkbuf_1 _4207_ (.A(_2145_),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _4208_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[90].S.IN1_L4 ),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _4209_ (.A(_2146_),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _4210_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[91].S.IN1_L4 ),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_1 _4211_ (.A(_2147_),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _4212_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[92].S.IN1_L4 ),
    .X(_2148_));
 sky130_fd_sc_hd__clkbuf_1 _4213_ (.A(_2148_),
    .X(_0601_));
 sky130_fd_sc_hd__and3_1 _4214_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[93].S.IN1_L4 ),
    .X(_2149_));
 sky130_fd_sc_hd__clkbuf_1 _4215_ (.A(_2149_),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _4216_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[94].S.IN1_L4 ),
    .X(_2150_));
 sky130_fd_sc_hd__clkbuf_1 _4217_ (.A(_2150_),
    .X(_0611_));
 sky130_fd_sc_hd__and3_1 _4218_ (.A(_2144_),
    .B(_2140_),
    .C(\stage_gen[1].mux_gen[95].S.IN1_L4 ),
    .X(_2151_));
 sky130_fd_sc_hd__clkbuf_1 _4219_ (.A(_2151_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _4220_ (.A(_2041_),
    .X(_2152_));
 sky130_fd_sc_hd__and3_1 _4221_ (.A(_2144_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[96].S.IN1_L4 ),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_1 _4222_ (.A(_2153_),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _4223_ (.A(_2144_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[97].S.IN1_L4 ),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _4224_ (.A(_2154_),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _4225_ (.A(_2144_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[98].S.IN1_L4 ),
    .X(_2155_));
 sky130_fd_sc_hd__clkbuf_1 _4226_ (.A(_2155_),
    .X(_0631_));
 sky130_fd_sc_hd__buf_2 _4227_ (.A(_2059_),
    .X(_2156_));
 sky130_fd_sc_hd__and3_1 _4228_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[99].S.IN1_L4 ),
    .X(_2157_));
 sky130_fd_sc_hd__clkbuf_1 _4229_ (.A(_2157_),
    .X(_0636_));
 sky130_fd_sc_hd__and3_1 _4230_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[100].S.IN1_L4 ),
    .X(_2158_));
 sky130_fd_sc_hd__clkbuf_1 _4231_ (.A(_2158_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _4232_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[101].S.IN1_L4 ),
    .X(_2159_));
 sky130_fd_sc_hd__clkbuf_1 _4233_ (.A(_2159_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_1 _4234_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[102].S.IN1_L4 ),
    .X(_2160_));
 sky130_fd_sc_hd__clkbuf_1 _4235_ (.A(_2160_),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _4236_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[103].S.IN1_L4 ),
    .X(_2161_));
 sky130_fd_sc_hd__clkbuf_1 _4237_ (.A(_2161_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _4238_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[104].S.IN1_L4 ),
    .X(_2162_));
 sky130_fd_sc_hd__clkbuf_1 _4239_ (.A(_2162_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_1 _4240_ (.A(_2156_),
    .B(_2152_),
    .C(\stage_gen[1].mux_gen[105].S.IN1_L4 ),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_1 _4241_ (.A(_2163_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_6 _4242_ (.A(_1360_),
    .X(_2164_));
 sky130_fd_sc_hd__clkbuf_4 _4243_ (.A(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__and3_1 _4244_ (.A(_2156_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[106].S.IN1_L4 ),
    .X(_2166_));
 sky130_fd_sc_hd__clkbuf_1 _4245_ (.A(_2166_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _4246_ (.A(_2156_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[107].S.IN1_L4 ),
    .X(_2167_));
 sky130_fd_sc_hd__clkbuf_1 _4247_ (.A(_2167_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _4248_ (.A(_2156_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[108].S.IN1_L4 ),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_1 _4249_ (.A(_2168_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_4 _4250_ (.A(_2059_),
    .X(_2169_));
 sky130_fd_sc_hd__and3_1 _4251_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[109].S.IN1_L4 ),
    .X(_2170_));
 sky130_fd_sc_hd__clkbuf_1 _4252_ (.A(_2170_),
    .X(_0056_));
 sky130_fd_sc_hd__and3_1 _4253_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[110].S.IN1_L4 ),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_1 _4254_ (.A(_2171_),
    .X(_0066_));
 sky130_fd_sc_hd__and3_1 _4255_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[111].S.IN1_L4 ),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _4256_ (.A(_2172_),
    .X(_0071_));
 sky130_fd_sc_hd__and3_1 _4257_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[112].S.IN1_L4 ),
    .X(_2173_));
 sky130_fd_sc_hd__clkbuf_1 _4258_ (.A(_2173_),
    .X(_0076_));
 sky130_fd_sc_hd__and3_1 _4259_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[113].S.IN1_L4 ),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _4260_ (.A(_2174_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _4261_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[114].S.IN1_L4 ),
    .X(_2175_));
 sky130_fd_sc_hd__clkbuf_1 _4262_ (.A(_2175_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _4263_ (.A(_2169_),
    .B(_2165_),
    .C(\stage_gen[1].mux_gen[115].S.IN1_L4 ),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _4264_ (.A(_2176_),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_4 _4265_ (.A(_2164_),
    .X(_2177_));
 sky130_fd_sc_hd__and3_1 _4266_ (.A(_2169_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[116].S.IN1_L4 ),
    .X(_2178_));
 sky130_fd_sc_hd__clkbuf_1 _4267_ (.A(_2178_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _4268_ (.A(_2169_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[117].S.IN1_L4 ),
    .X(_2179_));
 sky130_fd_sc_hd__clkbuf_1 _4269_ (.A(_2179_),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _4270_ (.A(_2169_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[118].S.IN1_L4 ),
    .X(_2180_));
 sky130_fd_sc_hd__clkbuf_1 _4271_ (.A(_2180_),
    .X(_0106_));
 sky130_fd_sc_hd__and3_1 _4272_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[119].S.IN1_L4 ),
    .X(_2181_));
 sky130_fd_sc_hd__clkbuf_1 _4273_ (.A(_2181_),
    .X(_0111_));
 sky130_fd_sc_hd__and3_1 _4274_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[120].S.IN1_L4 ),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_1 _4275_ (.A(_2182_),
    .X(_0121_));
 sky130_fd_sc_hd__and3_1 _4276_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[121].S.IN1_L4 ),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _4277_ (.A(_2183_),
    .X(_0126_));
 sky130_fd_sc_hd__and3_1 _4278_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[122].S.IN1_L4 ),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_1 _4279_ (.A(_2184_),
    .X(_0131_));
 sky130_fd_sc_hd__and3_1 _4280_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[123].S.IN1_L4 ),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _4281_ (.A(_2185_),
    .X(_0136_));
 sky130_fd_sc_hd__and3_1 _4282_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[124].S.IN1_L4 ),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _4283_ (.A(_2186_),
    .X(_0141_));
 sky130_fd_sc_hd__and3_1 _4284_ (.A(_2046_),
    .B(_2177_),
    .C(\stage_gen[1].mux_gen[125].S.IN1_L4 ),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_1 _4285_ (.A(_2187_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_4 _4286_ (.A(_2164_),
    .X(_2188_));
 sky130_fd_sc_hd__and3_1 _4287_ (.A(_2046_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[126].S.IN1_L4 ),
    .X(_2189_));
 sky130_fd_sc_hd__clkbuf_1 _4288_ (.A(_2189_),
    .X(_0151_));
 sky130_fd_sc_hd__and3_1 _4289_ (.A(_2046_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[127].S.IN1_L4 ),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_1 _4290_ (.A(_2190_),
    .X(_0156_));
 sky130_fd_sc_hd__and3_1 _4291_ (.A(_1513_),
    .B(_1965_),
    .C(\stage_gen[2].mux_gen[0].S.IN1_L4 ),
    .X(_2191_));
 sky130_fd_sc_hd__clkbuf_1 _4292_ (.A(_2191_),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _4293_ (.A(_1513_),
    .B(_1965_),
    .C(\stage_gen[2].mux_gen[1].S.IN1_L4 ),
    .X(_2192_));
 sky130_fd_sc_hd__clkbuf_1 _4294_ (.A(_2192_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_4 _4295_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .X(_2193_));
 sky130_fd_sc_hd__buf_2 _4296_ (.A(_1682_),
    .X(_2194_));
 sky130_fd_sc_hd__and3_1 _4297_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[2].S.IN1_L4 ),
    .X(_2195_));
 sky130_fd_sc_hd__clkbuf_1 _4298_ (.A(_2195_),
    .X(_0758_));
 sky130_fd_sc_hd__and3_1 _4299_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[3].S.IN1_L4 ),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _4300_ (.A(_2196_),
    .X(_0813_));
 sky130_fd_sc_hd__and3_1 _4301_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[4].S.IN1_L4 ),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _4302_ (.A(_2197_),
    .X(_0868_));
 sky130_fd_sc_hd__and3_1 _4303_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[5].S.IN1_L4 ),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _4304_ (.A(_2198_),
    .X(_0923_));
 sky130_fd_sc_hd__and3_1 _4305_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[6].S.IN1_L4 ),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _4306_ (.A(_2199_),
    .X(_0948_));
 sky130_fd_sc_hd__and3_1 _4307_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[7].S.IN1_L4 ),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _4308_ (.A(_2200_),
    .X(_0953_));
 sky130_fd_sc_hd__and3_1 _4309_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[8].S.IN1_L4 ),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_2201_),
    .X(_0958_));
 sky130_fd_sc_hd__and3_1 _4311_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[9].S.IN1_L4 ),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_1 _4312_ (.A(_2202_),
    .X(_0963_));
 sky130_fd_sc_hd__and3_1 _4313_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[10].S.IN1_L4 ),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_2203_),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _4315_ (.A(_2193_),
    .B(_2194_),
    .C(\stage_gen[2].mux_gen[11].S.IN1_L4 ),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _4316_ (.A(_2204_),
    .X(_0658_));
 sky130_fd_sc_hd__buf_2 _4317_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_2 _4318_ (.A(_1682_),
    .X(_2206_));
 sky130_fd_sc_hd__and3_1 _4319_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[12].S.IN1_L4 ),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_1 _4320_ (.A(_2207_),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _4321_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[13].S.IN1_L4 ),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_1 _4322_ (.A(_2208_),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _4323_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[14].S.IN1_L4 ),
    .X(_2209_));
 sky130_fd_sc_hd__clkbuf_1 _4324_ (.A(_2209_),
    .X(_0673_));
 sky130_fd_sc_hd__and3_1 _4325_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[15].S.IN1_L4 ),
    .X(_2210_));
 sky130_fd_sc_hd__clkbuf_1 _4326_ (.A(_2210_),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _4327_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[16].S.IN1_L4 ),
    .X(_2211_));
 sky130_fd_sc_hd__clkbuf_1 _4328_ (.A(_2211_),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _4329_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[17].S.IN1_L4 ),
    .X(_2212_));
 sky130_fd_sc_hd__clkbuf_1 _4330_ (.A(_2212_),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _4331_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[18].S.IN1_L4 ),
    .X(_2213_));
 sky130_fd_sc_hd__clkbuf_1 _4332_ (.A(_2213_),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _4333_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[19].S.IN1_L4 ),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_1 _4334_ (.A(_2214_),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _4335_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[20].S.IN1_L4 ),
    .X(_2215_));
 sky130_fd_sc_hd__clkbuf_1 _4336_ (.A(_2215_),
    .X(_0708_));
 sky130_fd_sc_hd__and3_1 _4337_ (.A(_2205_),
    .B(_2206_),
    .C(\stage_gen[2].mux_gen[21].S.IN1_L4 ),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_1 _4338_ (.A(_2216_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_2 _4339_ (.A(\stage_gen[2].genblk1.clks.clk_o ),
    .X(_2217_));
 sky130_fd_sc_hd__buf_2 _4340_ (.A(_1682_),
    .X(_2218_));
 sky130_fd_sc_hd__and3_1 _4341_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[22].S.IN1_L4 ),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _4342_ (.A(_2219_),
    .X(_0718_));
 sky130_fd_sc_hd__and3_1 _4343_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[23].S.IN1_L4 ),
    .X(_2220_));
 sky130_fd_sc_hd__clkbuf_1 _4344_ (.A(_2220_),
    .X(_0723_));
 sky130_fd_sc_hd__and3_1 _4345_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[24].S.IN1_L4 ),
    .X(_2221_));
 sky130_fd_sc_hd__clkbuf_1 _4346_ (.A(_2221_),
    .X(_0728_));
 sky130_fd_sc_hd__and3_1 _4347_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[25].S.IN1_L4 ),
    .X(_2222_));
 sky130_fd_sc_hd__clkbuf_1 _4348_ (.A(_2222_),
    .X(_0733_));
 sky130_fd_sc_hd__and3_1 _4349_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[26].S.IN1_L4 ),
    .X(_2223_));
 sky130_fd_sc_hd__clkbuf_1 _4350_ (.A(_2223_),
    .X(_0738_));
 sky130_fd_sc_hd__and3_1 _4351_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[27].S.IN1_L4 ),
    .X(_2224_));
 sky130_fd_sc_hd__clkbuf_1 _4352_ (.A(_2224_),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _4353_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[28].S.IN1_L4 ),
    .X(_2225_));
 sky130_fd_sc_hd__clkbuf_1 _4354_ (.A(_2225_),
    .X(_0748_));
 sky130_fd_sc_hd__and3_1 _4355_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[29].S.IN1_L4 ),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_1 _4356_ (.A(_2226_),
    .X(_0753_));
 sky130_fd_sc_hd__and3_1 _4357_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[30].S.IN1_L4 ),
    .X(_2227_));
 sky130_fd_sc_hd__clkbuf_1 _4358_ (.A(_2227_),
    .X(_0763_));
 sky130_fd_sc_hd__and3_1 _4359_ (.A(_2217_),
    .B(_2218_),
    .C(\stage_gen[2].mux_gen[31].S.IN1_L4 ),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_1 _4360_ (.A(_2228_),
    .X(_0768_));
 sky130_fd_sc_hd__and3_1 _4361_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[32].S.IN1_L4 ),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_1 _4362_ (.A(_2229_),
    .X(_0773_));
 sky130_fd_sc_hd__and3_1 _4363_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[33].S.IN1_L4 ),
    .X(_2230_));
 sky130_fd_sc_hd__clkbuf_1 _4364_ (.A(_2230_),
    .X(_0778_));
 sky130_fd_sc_hd__and3_1 _4365_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[34].S.IN1_L4 ),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_1 _4366_ (.A(_2231_),
    .X(_0783_));
 sky130_fd_sc_hd__and3_1 _4367_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[35].S.IN1_L4 ),
    .X(_2232_));
 sky130_fd_sc_hd__clkbuf_1 _4368_ (.A(_2232_),
    .X(_0788_));
 sky130_fd_sc_hd__and3_1 _4369_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[36].S.IN1_L4 ),
    .X(_2233_));
 sky130_fd_sc_hd__clkbuf_1 _4370_ (.A(_2233_),
    .X(_0793_));
 sky130_fd_sc_hd__and3_1 _4371_ (.A(_1363_),
    .B(_1801_),
    .C(\stage_gen[2].mux_gen[37].S.IN1_L4 ),
    .X(_2234_));
 sky130_fd_sc_hd__clkbuf_1 _4372_ (.A(_2234_),
    .X(_0798_));
 sky130_fd_sc_hd__clkinv_4 _4373_ (.A(_1361_),
    .Y(_2235_));
 sky130_fd_sc_hd__nor2_8 _4374_ (.A(clknet_1_1__leaf__2017_),
    .B(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__buf_6 _4375_ (.A(clknet_1_0__leaf__2236_),
    .X(_1290_));
 sky130_fd_sc_hd__nor2_2 _4376_ (.A(_2027_),
    .B(clknet_1_1__leaf__2022_),
    .Y(_1288_));
 sky130_fd_sc_hd__clkbuf_4 _4377_ (.A(_1368_),
    .X(_2237_));
 sky130_fd_sc_hd__buf_4 _4378_ (.A(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__buf_4 _4379_ (.A(_2032_),
    .X(_2239_));
 sky130_fd_sc_hd__a22o_1 _4380_ (.A1(_2238_),
    .A2(\stage_gen[1].mux_gen[0].S.IN1_L1 ),
    .B1(_2239_),
    .B2(net1),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _4381_ (.A(_1371_),
    .X(_2240_));
 sky130_fd_sc_hd__and3_1 _4382_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[0].S.IN1_L2 ),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_1 _4383_ (.A(_2241_),
    .X(_0002_));
 sky130_fd_sc_hd__a21o_1 _4384_ (.A1(\stage_gen[1].mux_gen[0].S.IN1_L1 ),
    .A2(net372),
    .B1(_0002_),
    .X(_0001_));
 sky130_fd_sc_hd__a21o_1 _4385_ (.A1(net112),
    .A2(net281),
    .B1(_0004_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_4 _4386_ (.A(_2033_),
    .X(_2242_));
 sky130_fd_sc_hd__buf_4 _4387_ (.A(_1373_),
    .X(_2243_));
 sky130_fd_sc_hd__buf_4 _4388_ (.A(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__a22o_1 _4389_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[1].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net179),
    .X(_0197_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[1].S.IN1_L2 ),
    .X(_2245_));
 sky130_fd_sc_hd__clkbuf_1 _4391_ (.A(_2245_),
    .X(_0199_));
 sky130_fd_sc_hd__a21o_1 _4392_ (.A1(\stage_gen[1].mux_gen[1].S.IN1_L1 ),
    .A2(net367),
    .B1(_0199_),
    .X(_0198_));
 sky130_fd_sc_hd__a21o_1 _4393_ (.A1(net190),
    .A2(net282),
    .B1(_0201_),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _4394_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[2].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net201),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _4395_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[2].S.IN1_L2 ),
    .X(_2246_));
 sky130_fd_sc_hd__clkbuf_1 _4396_ (.A(_2246_),
    .X(_0254_));
 sky130_fd_sc_hd__a21o_1 _4397_ (.A1(\stage_gen[1].mux_gen[2].S.IN1_L1 ),
    .A2(net367),
    .B1(_0254_),
    .X(_0253_));
 sky130_fd_sc_hd__a21o_1 _4398_ (.A1(net212),
    .A2(net276),
    .B1(_0256_),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _4399_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[3].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net223),
    .X(_0307_));
 sky130_fd_sc_hd__and3_1 _4400_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[3].S.IN1_L2 ),
    .X(_2247_));
 sky130_fd_sc_hd__clkbuf_1 _4401_ (.A(_2247_),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _4402_ (.A1(\stage_gen[1].mux_gen[3].S.IN1_L1 ),
    .A2(net366),
    .B1(_0309_),
    .X(_0308_));
 sky130_fd_sc_hd__a21o_1 _4403_ (.A1(net234),
    .A2(net280),
    .B1(_0311_),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _4404_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[4].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net245),
    .X(_0362_));
 sky130_fd_sc_hd__and3_1 _4405_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[4].S.IN1_L2 ),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_1 _4406_ (.A(_2248_),
    .X(_0364_));
 sky130_fd_sc_hd__a21o_1 _4407_ (.A1(\stage_gen[1].mux_gen[4].S.IN1_L1 ),
    .A2(net367),
    .B1(_0364_),
    .X(_0363_));
 sky130_fd_sc_hd__a21o_1 _4408_ (.A1(net256),
    .A2(net276),
    .B1(_0366_),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _4409_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[5].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net12),
    .X(_0417_));
 sky130_fd_sc_hd__and3_1 _4410_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[5].S.IN1_L2 ),
    .X(_2249_));
 sky130_fd_sc_hd__clkbuf_1 _4411_ (.A(_2249_),
    .X(_0419_));
 sky130_fd_sc_hd__a21o_1 _4412_ (.A1(\stage_gen[1].mux_gen[5].S.IN1_L1 ),
    .A2(net370),
    .B1(_0419_),
    .X(_0418_));
 sky130_fd_sc_hd__a21o_1 _4413_ (.A1(net23),
    .A2(net277),
    .B1(_0421_),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _4414_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[6].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net34),
    .X(_0472_));
 sky130_fd_sc_hd__and3_1 _4415_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[6].S.IN1_L2 ),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_1 _4416_ (.A(_2250_),
    .X(_0474_));
 sky130_fd_sc_hd__a21o_1 _4417_ (.A1(\stage_gen[1].mux_gen[6].S.IN1_L1 ),
    .A2(net360),
    .B1(_0474_),
    .X(_0473_));
 sky130_fd_sc_hd__a21o_1 _4418_ (.A1(net45),
    .A2(net274),
    .B1(_0476_),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _4419_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[7].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net56),
    .X(_0527_));
 sky130_fd_sc_hd__and3_1 _4420_ (.A(_2240_),
    .B(_2188_),
    .C(\stage_gen[1].mux_gen[7].S.IN1_L2 ),
    .X(_2251_));
 sky130_fd_sc_hd__clkbuf_1 _4421_ (.A(_2251_),
    .X(_0529_));
 sky130_fd_sc_hd__a21o_1 _4422_ (.A1(\stage_gen[1].mux_gen[7].S.IN1_L1 ),
    .A2(net369),
    .B1(_0529_),
    .X(_0528_));
 sky130_fd_sc_hd__a21o_1 _4423_ (.A1(net67),
    .A2(net277),
    .B1(_0531_),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _4424_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[8].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net78),
    .X(_0582_));
 sky130_fd_sc_hd__buf_2 _4425_ (.A(_2164_),
    .X(_2252_));
 sky130_fd_sc_hd__and3_1 _4426_ (.A(_2240_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[8].S.IN1_L2 ),
    .X(_2253_));
 sky130_fd_sc_hd__clkbuf_1 _4427_ (.A(_2253_),
    .X(_0584_));
 sky130_fd_sc_hd__a21o_1 _4428_ (.A1(\stage_gen[1].mux_gen[8].S.IN1_L1 ),
    .A2(net335),
    .B1(_0584_),
    .X(_0583_));
 sky130_fd_sc_hd__a21o_1 _4429_ (.A1(net89),
    .A2(net278),
    .B1(_0586_),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _4430_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[9].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net100),
    .X(_0637_));
 sky130_fd_sc_hd__buf_4 _4431_ (.A(_1368_),
    .X(_2254_));
 sky130_fd_sc_hd__clkbuf_4 _4432_ (.A(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__clkbuf_4 _4433_ (.A(_1371_),
    .X(_2256_));
 sky130_fd_sc_hd__buf_2 _4434_ (.A(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__and3_1 _4435_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[9].S.IN1_L2 ),
    .X(_2258_));
 sky130_fd_sc_hd__clkbuf_1 _4436_ (.A(_2258_),
    .X(_0639_));
 sky130_fd_sc_hd__a21o_1 _4437_ (.A1(\stage_gen[1].mux_gen[9].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0639_),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_4 _4438_ (.A(_1373_),
    .X(_2259_));
 sky130_fd_sc_hd__clkbuf_4 _4439_ (.A(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a21o_1 _4440_ (.A1(net111),
    .A2(_2260_),
    .B1(_0641_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _4441_ (.A1(_2242_),
    .A2(\stage_gen[1].mux_gen[10].S.IN1_L1 ),
    .B1(_2244_),
    .B2(net123),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _4442_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[10].S.IN1_L2 ),
    .X(_2261_));
 sky130_fd_sc_hd__clkbuf_1 _4443_ (.A(_2261_),
    .X(_0059_));
 sky130_fd_sc_hd__a21o_1 _4444_ (.A1(\stage_gen[1].mux_gen[10].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0059_),
    .X(_0058_));
 sky130_fd_sc_hd__a21o_1 _4445_ (.A1(net134),
    .A2(_2260_),
    .B1(_0061_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_4 _4446_ (.A(_2033_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_4 _4447_ (.A(_2243_),
    .X(_2263_));
 sky130_fd_sc_hd__a22o_1 _4448_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[11].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net145),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _4449_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[11].S.IN1_L2 ),
    .X(_2264_));
 sky130_fd_sc_hd__clkbuf_1 _4450_ (.A(_2264_),
    .X(_0114_));
 sky130_fd_sc_hd__a21o_1 _4451_ (.A1(\stage_gen[1].mux_gen[11].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0114_),
    .X(_0113_));
 sky130_fd_sc_hd__a21o_1 _4452_ (.A1(net156),
    .A2(_2260_),
    .B1(_0116_),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _4453_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[12].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net167),
    .X(_0157_));
 sky130_fd_sc_hd__and3_1 _4454_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[12].S.IN1_L2 ),
    .X(_2265_));
 sky130_fd_sc_hd__clkbuf_1 _4455_ (.A(_2265_),
    .X(_0159_));
 sky130_fd_sc_hd__a21o_1 _4456_ (.A1(\stage_gen[1].mux_gen[12].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0159_),
    .X(_0158_));
 sky130_fd_sc_hd__a21o_1 _4457_ (.A1(net174),
    .A2(_2260_),
    .B1(_0161_),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _4458_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[13].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net175),
    .X(_0162_));
 sky130_fd_sc_hd__and3_1 _4459_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[13].S.IN1_L2 ),
    .X(_2266_));
 sky130_fd_sc_hd__clkbuf_1 _4460_ (.A(_2266_),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_1 _4461_ (.A1(\stage_gen[1].mux_gen[13].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0164_),
    .X(_0163_));
 sky130_fd_sc_hd__a21o_1 _4462_ (.A1(net176),
    .A2(_2260_),
    .B1(_0166_),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _4463_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[14].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net177),
    .X(_0167_));
 sky130_fd_sc_hd__and3_1 _4464_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[14].S.IN1_L2 ),
    .X(_2267_));
 sky130_fd_sc_hd__clkbuf_1 _4465_ (.A(_2267_),
    .X(_0169_));
 sky130_fd_sc_hd__a21o_1 _4466_ (.A1(\stage_gen[1].mux_gen[14].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0169_),
    .X(_0168_));
 sky130_fd_sc_hd__a21o_1 _4467_ (.A1(net178),
    .A2(_2260_),
    .B1(_0171_),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _4468_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[15].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net180),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _4469_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[15].S.IN1_L2 ),
    .X(_2268_));
 sky130_fd_sc_hd__clkbuf_1 _4470_ (.A(_2268_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _4471_ (.A1(\stage_gen[1].mux_gen[15].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0174_),
    .X(_0173_));
 sky130_fd_sc_hd__a21o_1 _4472_ (.A1(net181),
    .A2(_2260_),
    .B1(_0176_),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _4473_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[16].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net182),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _4474_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[16].S.IN1_L2 ),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_1 _4475_ (.A(_2269_),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_1 _4476_ (.A1(\stage_gen[1].mux_gen[16].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0179_),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_1 _4477_ (.A1(net183),
    .A2(_2260_),
    .B1(_0181_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _4478_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[17].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net184),
    .X(_0182_));
 sky130_fd_sc_hd__and3_1 _4479_ (.A(_2257_),
    .B(_2252_),
    .C(\stage_gen[1].mux_gen[17].S.IN1_L2 ),
    .X(_2270_));
 sky130_fd_sc_hd__clkbuf_1 _4480_ (.A(_2270_),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _4481_ (.A1(\stage_gen[1].mux_gen[17].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0184_),
    .X(_0183_));
 sky130_fd_sc_hd__a21o_1 _4482_ (.A1(net185),
    .A2(_2260_),
    .B1(_0186_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _4483_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[18].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net186),
    .X(_0187_));
 sky130_fd_sc_hd__buf_2 _4484_ (.A(_2164_),
    .X(_2271_));
 sky130_fd_sc_hd__and3_1 _4485_ (.A(_2257_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[18].S.IN1_L2 ),
    .X(_2272_));
 sky130_fd_sc_hd__clkbuf_1 _4486_ (.A(_2272_),
    .X(_0189_));
 sky130_fd_sc_hd__a21o_1 _4487_ (.A1(\stage_gen[1].mux_gen[18].S.IN1_L1 ),
    .A2(_2255_),
    .B1(_0189_),
    .X(_0188_));
 sky130_fd_sc_hd__a21o_1 _4488_ (.A1(net187),
    .A2(_2260_),
    .B1(_0191_),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_1 _4489_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[19].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net188),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _4490_ (.A(_2254_),
    .X(_2273_));
 sky130_fd_sc_hd__buf_4 _4491_ (.A(_1371_),
    .X(_2274_));
 sky130_fd_sc_hd__clkbuf_2 _4492_ (.A(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__and3_1 _4493_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[19].S.IN1_L2 ),
    .X(_2276_));
 sky130_fd_sc_hd__clkbuf_1 _4494_ (.A(_2276_),
    .X(_0194_));
 sky130_fd_sc_hd__a21o_1 _4495_ (.A1(\stage_gen[1].mux_gen[19].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0194_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_4 _4496_ (.A(_2259_),
    .X(_2277_));
 sky130_fd_sc_hd__a21o_1 _4497_ (.A1(net189),
    .A2(_2277_),
    .B1(_0196_),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _4498_ (.A1(_2262_),
    .A2(\stage_gen[1].mux_gen[20].S.IN1_L1 ),
    .B1(_2263_),
    .B2(net191),
    .X(_0202_));
 sky130_fd_sc_hd__and3_1 _4499_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[20].S.IN1_L2 ),
    .X(_2278_));
 sky130_fd_sc_hd__clkbuf_1 _4500_ (.A(_2278_),
    .X(_0204_));
 sky130_fd_sc_hd__a21o_1 _4501_ (.A1(\stage_gen[1].mux_gen[20].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0204_),
    .X(_0203_));
 sky130_fd_sc_hd__a21o_1 _4502_ (.A1(net192),
    .A2(_2277_),
    .B1(_0206_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_4 _4503_ (.A(_2033_),
    .X(_2279_));
 sky130_fd_sc_hd__buf_2 _4504_ (.A(_2243_),
    .X(_2280_));
 sky130_fd_sc_hd__a22o_1 _4505_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[21].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net193),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _4506_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[21].S.IN1_L2 ),
    .X(_2281_));
 sky130_fd_sc_hd__clkbuf_1 _4507_ (.A(_2281_),
    .X(_0209_));
 sky130_fd_sc_hd__a21o_1 _4508_ (.A1(\stage_gen[1].mux_gen[21].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0209_),
    .X(_0208_));
 sky130_fd_sc_hd__a21o_1 _4509_ (.A1(net194),
    .A2(_2277_),
    .B1(_0211_),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _4510_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[22].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net195),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _4511_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[22].S.IN1_L2 ),
    .X(_2282_));
 sky130_fd_sc_hd__clkbuf_1 _4512_ (.A(_2282_),
    .X(_0214_));
 sky130_fd_sc_hd__a21o_1 _4513_ (.A1(\stage_gen[1].mux_gen[22].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0214_),
    .X(_0213_));
 sky130_fd_sc_hd__a21o_1 _4514_ (.A1(net196),
    .A2(_2277_),
    .B1(_0216_),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _4515_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[23].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net197),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _4516_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[23].S.IN1_L2 ),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _4517_ (.A(_2283_),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _4518_ (.A1(\stage_gen[1].mux_gen[23].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0219_),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _4519_ (.A1(net198),
    .A2(_2277_),
    .B1(_0221_),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _4520_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[24].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net199),
    .X(_0222_));
 sky130_fd_sc_hd__and3_1 _4521_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[24].S.IN1_L2 ),
    .X(_2284_));
 sky130_fd_sc_hd__clkbuf_1 _4522_ (.A(_2284_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _4523_ (.A1(\stage_gen[1].mux_gen[24].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0224_),
    .X(_0223_));
 sky130_fd_sc_hd__a21o_1 _4524_ (.A1(net200),
    .A2(_2277_),
    .B1(_0226_),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _4525_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[25].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net202),
    .X(_0227_));
 sky130_fd_sc_hd__and3_1 _4526_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[25].S.IN1_L2 ),
    .X(_2285_));
 sky130_fd_sc_hd__clkbuf_1 _4527_ (.A(_2285_),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_1 _4528_ (.A1(\stage_gen[1].mux_gen[25].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0229_),
    .X(_0228_));
 sky130_fd_sc_hd__a21o_1 _4529_ (.A1(net203),
    .A2(_2277_),
    .B1(_0231_),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _4530_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[26].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net204),
    .X(_0232_));
 sky130_fd_sc_hd__and3_1 _4531_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[26].S.IN1_L2 ),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _4532_ (.A(_2286_),
    .X(_0234_));
 sky130_fd_sc_hd__a21o_1 _4533_ (.A1(\stage_gen[1].mux_gen[26].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0234_),
    .X(_0233_));
 sky130_fd_sc_hd__a21o_1 _4534_ (.A1(net205),
    .A2(_2277_),
    .B1(_0236_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _4535_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[27].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net206),
    .X(_0237_));
 sky130_fd_sc_hd__and3_1 _4536_ (.A(_2275_),
    .B(_2271_),
    .C(\stage_gen[1].mux_gen[27].S.IN1_L2 ),
    .X(_2287_));
 sky130_fd_sc_hd__clkbuf_1 _4537_ (.A(_2287_),
    .X(_0239_));
 sky130_fd_sc_hd__a21o_1 _4538_ (.A1(\stage_gen[1].mux_gen[27].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0239_),
    .X(_0238_));
 sky130_fd_sc_hd__a21o_1 _4539_ (.A1(net207),
    .A2(_2277_),
    .B1(_0241_),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _4540_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[28].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net208),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_2 _4541_ (.A(_2164_),
    .X(_2288_));
 sky130_fd_sc_hd__and3_1 _4542_ (.A(_2275_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[28].S.IN1_L2 ),
    .X(_2289_));
 sky130_fd_sc_hd__clkbuf_1 _4543_ (.A(_2289_),
    .X(_0244_));
 sky130_fd_sc_hd__a21o_1 _4544_ (.A1(\stage_gen[1].mux_gen[28].S.IN1_L1 ),
    .A2(_2273_),
    .B1(_0244_),
    .X(_0243_));
 sky130_fd_sc_hd__a21o_1 _4545_ (.A1(net209),
    .A2(_2277_),
    .B1(_0246_),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _4546_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[29].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net210),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_4 _4547_ (.A(_2254_),
    .X(_2290_));
 sky130_fd_sc_hd__clkbuf_2 _4548_ (.A(_2274_),
    .X(_2291_));
 sky130_fd_sc_hd__and3_1 _4549_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[29].S.IN1_L2 ),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _4550_ (.A(_2292_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _4551_ (.A1(\stage_gen[1].mux_gen[29].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0249_),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_4 _4552_ (.A(_2259_),
    .X(_2293_));
 sky130_fd_sc_hd__a21o_1 _4553_ (.A1(net211),
    .A2(_2293_),
    .B1(_0251_),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _4554_ (.A1(_2279_),
    .A2(\stage_gen[1].mux_gen[30].S.IN1_L1 ),
    .B1(_2280_),
    .B2(net213),
    .X(_0257_));
 sky130_fd_sc_hd__and3_1 _4555_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[30].S.IN1_L2 ),
    .X(_2294_));
 sky130_fd_sc_hd__clkbuf_1 _4556_ (.A(_2294_),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _4557_ (.A1(\stage_gen[1].mux_gen[30].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0259_),
    .X(_0258_));
 sky130_fd_sc_hd__a21o_1 _4558_ (.A1(net214),
    .A2(_2293_),
    .B1(_0261_),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_4 _4559_ (.A(_2237_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_4 _4560_ (.A(_2243_),
    .X(_2296_));
 sky130_fd_sc_hd__a22o_1 _4561_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[31].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net215),
    .X(_0262_));
 sky130_fd_sc_hd__and3_1 _4562_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[31].S.IN1_L2 ),
    .X(_2297_));
 sky130_fd_sc_hd__clkbuf_1 _4563_ (.A(_2297_),
    .X(_0264_));
 sky130_fd_sc_hd__a21o_1 _4564_ (.A1(\stage_gen[1].mux_gen[31].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0264_),
    .X(_0263_));
 sky130_fd_sc_hd__a21o_1 _4565_ (.A1(net216),
    .A2(_2293_),
    .B1(_0266_),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _4566_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[32].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net217),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _4567_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[32].S.IN1_L2 ),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _4568_ (.A(_2298_),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_1 _4569_ (.A1(\stage_gen[1].mux_gen[32].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0269_),
    .X(_0268_));
 sky130_fd_sc_hd__a21o_1 _4570_ (.A1(net218),
    .A2(_2293_),
    .B1(_0271_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _4571_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[33].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net219),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _4572_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[33].S.IN1_L2 ),
    .X(_2299_));
 sky130_fd_sc_hd__clkbuf_1 _4573_ (.A(_2299_),
    .X(_0274_));
 sky130_fd_sc_hd__a21o_1 _4574_ (.A1(\stage_gen[1].mux_gen[33].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0274_),
    .X(_0273_));
 sky130_fd_sc_hd__a21o_1 _4575_ (.A1(net220),
    .A2(_2293_),
    .B1(_0276_),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[34].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net221),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _4577_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[34].S.IN1_L2 ),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_1 _4578_ (.A(_2300_),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _4579_ (.A1(\stage_gen[1].mux_gen[34].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0279_),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _4580_ (.A1(net222),
    .A2(_2293_),
    .B1(_0281_),
    .X(_0280_));
 sky130_fd_sc_hd__a22o_1 _4581_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[35].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net224),
    .X(_0282_));
 sky130_fd_sc_hd__and3_1 _4582_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[35].S.IN1_L2 ),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _4583_ (.A(_2301_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_1 _4584_ (.A1(\stage_gen[1].mux_gen[35].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0284_),
    .X(_0283_));
 sky130_fd_sc_hd__a21o_1 _4585_ (.A1(net225),
    .A2(_2293_),
    .B1(_0286_),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[36].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net226),
    .X(_0287_));
 sky130_fd_sc_hd__and3_1 _4587_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[36].S.IN1_L2 ),
    .X(_2302_));
 sky130_fd_sc_hd__clkbuf_1 _4588_ (.A(_2302_),
    .X(_0289_));
 sky130_fd_sc_hd__a21o_1 _4589_ (.A1(\stage_gen[1].mux_gen[36].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0289_),
    .X(_0288_));
 sky130_fd_sc_hd__a21o_1 _4590_ (.A1(net227),
    .A2(_2293_),
    .B1(_0291_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _4591_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[37].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net228),
    .X(_0292_));
 sky130_fd_sc_hd__and3_1 _4592_ (.A(_2291_),
    .B(_2288_),
    .C(\stage_gen[1].mux_gen[37].S.IN1_L2 ),
    .X(_2303_));
 sky130_fd_sc_hd__clkbuf_1 _4593_ (.A(_2303_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _4594_ (.A1(\stage_gen[1].mux_gen[37].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0294_),
    .X(_0293_));
 sky130_fd_sc_hd__a21o_1 _4595_ (.A1(net229),
    .A2(_2293_),
    .B1(_0296_),
    .X(_0295_));
 sky130_fd_sc_hd__a22o_1 _4596_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[38].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net230),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _4597_ (.A(_2164_),
    .X(_2304_));
 sky130_fd_sc_hd__and3_1 _4598_ (.A(_2291_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[38].S.IN1_L2 ),
    .X(_2305_));
 sky130_fd_sc_hd__clkbuf_1 _4599_ (.A(_2305_),
    .X(_0299_));
 sky130_fd_sc_hd__a21o_1 _4600_ (.A1(\stage_gen[1].mux_gen[38].S.IN1_L1 ),
    .A2(_2290_),
    .B1(_0299_),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_1 _4601_ (.A1(net231),
    .A2(_2293_),
    .B1(_0301_),
    .X(_0300_));
 sky130_fd_sc_hd__a22o_1 _4602_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[39].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net232),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_4 _4603_ (.A(_2254_),
    .X(_2306_));
 sky130_fd_sc_hd__clkbuf_2 _4604_ (.A(_2274_),
    .X(_2307_));
 sky130_fd_sc_hd__and3_1 _4605_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[39].S.IN1_L2 ),
    .X(_2308_));
 sky130_fd_sc_hd__clkbuf_1 _4606_ (.A(_2308_),
    .X(_0304_));
 sky130_fd_sc_hd__a21o_1 _4607_ (.A1(\stage_gen[1].mux_gen[39].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0304_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _4608_ (.A(_2032_),
    .X(_2309_));
 sky130_fd_sc_hd__a21o_1 _4609_ (.A1(net233),
    .A2(_2309_),
    .B1(_0306_),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _4610_ (.A1(_2295_),
    .A2(\stage_gen[1].mux_gen[40].S.IN1_L1 ),
    .B1(_2296_),
    .B2(net235),
    .X(_0312_));
 sky130_fd_sc_hd__and3_1 _4611_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[40].S.IN1_L2 ),
    .X(_2310_));
 sky130_fd_sc_hd__clkbuf_1 _4612_ (.A(_2310_),
    .X(_0314_));
 sky130_fd_sc_hd__a21o_1 _4613_ (.A1(\stage_gen[1].mux_gen[40].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0314_),
    .X(_0313_));
 sky130_fd_sc_hd__a21o_1 _4614_ (.A1(net236),
    .A2(_2309_),
    .B1(_0316_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_4 _4615_ (.A(_2237_),
    .X(_2311_));
 sky130_fd_sc_hd__clkbuf_4 _4616_ (.A(_2243_),
    .X(_2312_));
 sky130_fd_sc_hd__a22o_1 _4617_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[41].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net237),
    .X(_0317_));
 sky130_fd_sc_hd__and3_1 _4618_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[41].S.IN1_L2 ),
    .X(_2313_));
 sky130_fd_sc_hd__clkbuf_1 _4619_ (.A(_2313_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(\stage_gen[1].mux_gen[41].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0319_),
    .X(_0318_));
 sky130_fd_sc_hd__a21o_1 _4621_ (.A1(net238),
    .A2(_2309_),
    .B1(_0321_),
    .X(_0320_));
 sky130_fd_sc_hd__a22o_1 _4622_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[42].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net239),
    .X(_0322_));
 sky130_fd_sc_hd__and3_1 _4623_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[42].S.IN1_L2 ),
    .X(_2314_));
 sky130_fd_sc_hd__clkbuf_1 _4624_ (.A(_2314_),
    .X(_0324_));
 sky130_fd_sc_hd__a21o_1 _4625_ (.A1(\stage_gen[1].mux_gen[42].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0324_),
    .X(_0323_));
 sky130_fd_sc_hd__a21o_1 _4626_ (.A1(net240),
    .A2(_2309_),
    .B1(_0326_),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _4627_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[43].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net241),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _4628_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[43].S.IN1_L2 ),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_1 _4629_ (.A(_2315_),
    .X(_0329_));
 sky130_fd_sc_hd__a21o_1 _4630_ (.A1(\stage_gen[1].mux_gen[43].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0329_),
    .X(_0328_));
 sky130_fd_sc_hd__a21o_1 _4631_ (.A1(net242),
    .A2(_2309_),
    .B1(_0331_),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _4632_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[44].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net243),
    .X(_0332_));
 sky130_fd_sc_hd__and3_1 _4633_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[44].S.IN1_L2 ),
    .X(_2316_));
 sky130_fd_sc_hd__clkbuf_1 _4634_ (.A(_2316_),
    .X(_0334_));
 sky130_fd_sc_hd__a21o_1 _4635_ (.A1(\stage_gen[1].mux_gen[44].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0334_),
    .X(_0333_));
 sky130_fd_sc_hd__a21o_1 _4636_ (.A1(net244),
    .A2(_2309_),
    .B1(_0336_),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _4637_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[45].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net246),
    .X(_0337_));
 sky130_fd_sc_hd__and3_1 _4638_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[45].S.IN1_L2 ),
    .X(_2317_));
 sky130_fd_sc_hd__clkbuf_1 _4639_ (.A(_2317_),
    .X(_0339_));
 sky130_fd_sc_hd__a21o_1 _4640_ (.A1(\stage_gen[1].mux_gen[45].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0339_),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _4641_ (.A1(net247),
    .A2(_2309_),
    .B1(_0341_),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _4642_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[46].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net248),
    .X(_0342_));
 sky130_fd_sc_hd__and3_1 _4643_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[46].S.IN1_L2 ),
    .X(_2318_));
 sky130_fd_sc_hd__clkbuf_1 _4644_ (.A(_2318_),
    .X(_0344_));
 sky130_fd_sc_hd__a21o_1 _4645_ (.A1(\stage_gen[1].mux_gen[46].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0344_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _4646_ (.A1(net249),
    .A2(_2309_),
    .B1(_0346_),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _4647_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[47].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net250),
    .X(_0347_));
 sky130_fd_sc_hd__and3_1 _4648_ (.A(_2307_),
    .B(_2304_),
    .C(\stage_gen[1].mux_gen[47].S.IN1_L2 ),
    .X(_2319_));
 sky130_fd_sc_hd__clkbuf_1 _4649_ (.A(_2319_),
    .X(_0349_));
 sky130_fd_sc_hd__a21o_1 _4650_ (.A1(\stage_gen[1].mux_gen[47].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0349_),
    .X(_0348_));
 sky130_fd_sc_hd__a21o_1 _4651_ (.A1(net251),
    .A2(_2309_),
    .B1(_0351_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _4652_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[48].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net252),
    .X(_0352_));
 sky130_fd_sc_hd__buf_2 _4653_ (.A(_2164_),
    .X(_2320_));
 sky130_fd_sc_hd__and3_1 _4654_ (.A(_2307_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[48].S.IN1_L2 ),
    .X(_2321_));
 sky130_fd_sc_hd__clkbuf_1 _4655_ (.A(_2321_),
    .X(_0354_));
 sky130_fd_sc_hd__a21o_1 _4656_ (.A1(\stage_gen[1].mux_gen[48].S.IN1_L1 ),
    .A2(_2306_),
    .B1(_0354_),
    .X(_0353_));
 sky130_fd_sc_hd__a21o_1 _4657_ (.A1(net253),
    .A2(_2309_),
    .B1(_0356_),
    .X(_0355_));
 sky130_fd_sc_hd__a22o_1 _4658_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[49].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net254),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_4 _4659_ (.A(_2254_),
    .X(_2322_));
 sky130_fd_sc_hd__buf_2 _4660_ (.A(_2274_),
    .X(_2323_));
 sky130_fd_sc_hd__and3_1 _4661_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[49].S.IN1_L2 ),
    .X(_2324_));
 sky130_fd_sc_hd__clkbuf_1 _4662_ (.A(_2324_),
    .X(_0359_));
 sky130_fd_sc_hd__a21o_1 _4663_ (.A1(\stage_gen[1].mux_gen[49].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0359_),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_4 _4664_ (.A(_2032_),
    .X(_2325_));
 sky130_fd_sc_hd__a21o_1 _4665_ (.A1(net255),
    .A2(_2325_),
    .B1(_0361_),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _4666_ (.A1(_2311_),
    .A2(\stage_gen[1].mux_gen[50].S.IN1_L1 ),
    .B1(_2312_),
    .B2(net2),
    .X(_0367_));
 sky130_fd_sc_hd__and3_1 _4667_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[50].S.IN1_L2 ),
    .X(_2326_));
 sky130_fd_sc_hd__clkbuf_1 _4668_ (.A(_2326_),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _4669_ (.A1(\stage_gen[1].mux_gen[50].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0369_),
    .X(_0368_));
 sky130_fd_sc_hd__a21o_1 _4670_ (.A1(net3),
    .A2(_2325_),
    .B1(_0371_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_4 _4671_ (.A(_2237_),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_4 _4672_ (.A(_2259_),
    .X(_2328_));
 sky130_fd_sc_hd__a22o_1 _4673_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[51].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net4),
    .X(_0372_));
 sky130_fd_sc_hd__and3_1 _4674_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[51].S.IN1_L2 ),
    .X(_2329_));
 sky130_fd_sc_hd__clkbuf_1 _4675_ (.A(_2329_),
    .X(_0374_));
 sky130_fd_sc_hd__a21o_1 _4676_ (.A1(\stage_gen[1].mux_gen[51].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0374_),
    .X(_0373_));
 sky130_fd_sc_hd__a21o_1 _4677_ (.A1(net5),
    .A2(_2325_),
    .B1(_0376_),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _4678_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[52].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net6),
    .X(_0377_));
 sky130_fd_sc_hd__and3_1 _4679_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[52].S.IN1_L2 ),
    .X(_2330_));
 sky130_fd_sc_hd__clkbuf_1 _4680_ (.A(_2330_),
    .X(_0379_));
 sky130_fd_sc_hd__a21o_1 _4681_ (.A1(\stage_gen[1].mux_gen[52].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0379_),
    .X(_0378_));
 sky130_fd_sc_hd__a21o_1 _4682_ (.A1(net7),
    .A2(_2325_),
    .B1(_0381_),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _4683_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[53].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net8),
    .X(_0382_));
 sky130_fd_sc_hd__and3_1 _4684_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[53].S.IN1_L2 ),
    .X(_2331_));
 sky130_fd_sc_hd__clkbuf_1 _4685_ (.A(_2331_),
    .X(_0384_));
 sky130_fd_sc_hd__a21o_1 _4686_ (.A1(\stage_gen[1].mux_gen[53].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0384_),
    .X(_0383_));
 sky130_fd_sc_hd__a21o_1 _4687_ (.A1(net9),
    .A2(_2325_),
    .B1(_0386_),
    .X(_0385_));
 sky130_fd_sc_hd__a22o_1 _4688_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[54].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net10),
    .X(_0387_));
 sky130_fd_sc_hd__and3_1 _4689_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[54].S.IN1_L2 ),
    .X(_2332_));
 sky130_fd_sc_hd__clkbuf_1 _4690_ (.A(_2332_),
    .X(_0389_));
 sky130_fd_sc_hd__a21o_1 _4691_ (.A1(\stage_gen[1].mux_gen[54].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0389_),
    .X(_0388_));
 sky130_fd_sc_hd__a21o_1 _4692_ (.A1(net11),
    .A2(_2325_),
    .B1(_0391_),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _4693_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[55].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net13),
    .X(_0392_));
 sky130_fd_sc_hd__and3_1 _4694_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[55].S.IN1_L2 ),
    .X(_2333_));
 sky130_fd_sc_hd__clkbuf_1 _4695_ (.A(_2333_),
    .X(_0394_));
 sky130_fd_sc_hd__a21o_1 _4696_ (.A1(\stage_gen[1].mux_gen[55].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0394_),
    .X(_0393_));
 sky130_fd_sc_hd__a21o_1 _4697_ (.A1(net14),
    .A2(_2325_),
    .B1(_0396_),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _4698_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[56].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net15),
    .X(_0397_));
 sky130_fd_sc_hd__and3_1 _4699_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[56].S.IN1_L2 ),
    .X(_2334_));
 sky130_fd_sc_hd__clkbuf_1 _4700_ (.A(_2334_),
    .X(_0399_));
 sky130_fd_sc_hd__a21o_1 _4701_ (.A1(\stage_gen[1].mux_gen[56].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0399_),
    .X(_0398_));
 sky130_fd_sc_hd__a21o_1 _4702_ (.A1(net16),
    .A2(_2325_),
    .B1(_0401_),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_1 _4703_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[57].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net17),
    .X(_0402_));
 sky130_fd_sc_hd__and3_1 _4704_ (.A(_2323_),
    .B(_2320_),
    .C(\stage_gen[1].mux_gen[57].S.IN1_L2 ),
    .X(_2335_));
 sky130_fd_sc_hd__clkbuf_1 _4705_ (.A(_2335_),
    .X(_0404_));
 sky130_fd_sc_hd__a21o_1 _4706_ (.A1(\stage_gen[1].mux_gen[57].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0404_),
    .X(_0403_));
 sky130_fd_sc_hd__a21o_1 _4707_ (.A1(net18),
    .A2(_2325_),
    .B1(_0406_),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _4708_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[58].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net19),
    .X(_0407_));
 sky130_fd_sc_hd__buf_2 _4709_ (.A(_2164_),
    .X(_2336_));
 sky130_fd_sc_hd__and3_1 _4710_ (.A(_2323_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[58].S.IN1_L2 ),
    .X(_2337_));
 sky130_fd_sc_hd__clkbuf_1 _4711_ (.A(_2337_),
    .X(_0409_));
 sky130_fd_sc_hd__a21o_1 _4712_ (.A1(\stage_gen[1].mux_gen[58].S.IN1_L1 ),
    .A2(_2322_),
    .B1(_0409_),
    .X(_0408_));
 sky130_fd_sc_hd__a21o_1 _4713_ (.A1(net20),
    .A2(_2325_),
    .B1(_0411_),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _4714_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[59].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net21),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_4 _4715_ (.A(_2033_),
    .X(_2338_));
 sky130_fd_sc_hd__buf_2 _4716_ (.A(_2274_),
    .X(_2339_));
 sky130_fd_sc_hd__and3_1 _4717_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[59].S.IN1_L2 ),
    .X(_2340_));
 sky130_fd_sc_hd__clkbuf_1 _4718_ (.A(_2340_),
    .X(_0414_));
 sky130_fd_sc_hd__a21o_1 _4719_ (.A1(\stage_gen[1].mux_gen[59].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0414_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_4 _4720_ (.A(_2032_),
    .X(_2341_));
 sky130_fd_sc_hd__a21o_1 _4721_ (.A1(net22),
    .A2(_2341_),
    .B1(_0416_),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _4722_ (.A1(_2327_),
    .A2(\stage_gen[1].mux_gen[60].S.IN1_L1 ),
    .B1(_2328_),
    .B2(net24),
    .X(_0422_));
 sky130_fd_sc_hd__and3_1 _4723_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[60].S.IN1_L2 ),
    .X(_2342_));
 sky130_fd_sc_hd__clkbuf_1 _4724_ (.A(_2342_),
    .X(_0424_));
 sky130_fd_sc_hd__a21o_1 _4725_ (.A1(\stage_gen[1].mux_gen[60].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0424_),
    .X(_0423_));
 sky130_fd_sc_hd__a21o_1 _4726_ (.A1(net25),
    .A2(_2341_),
    .B1(_0426_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_4 _4727_ (.A(_2237_),
    .X(_2343_));
 sky130_fd_sc_hd__clkbuf_4 _4728_ (.A(_2259_),
    .X(_2344_));
 sky130_fd_sc_hd__a22o_1 _4729_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[61].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net26),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _4730_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[61].S.IN1_L2 ),
    .X(_2345_));
 sky130_fd_sc_hd__clkbuf_1 _4731_ (.A(_2345_),
    .X(_0429_));
 sky130_fd_sc_hd__a21o_1 _4732_ (.A1(\stage_gen[1].mux_gen[61].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0429_),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _4733_ (.A1(net27),
    .A2(_2341_),
    .B1(_0431_),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _4734_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[62].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net28),
    .X(_0432_));
 sky130_fd_sc_hd__and3_1 _4735_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[62].S.IN1_L2 ),
    .X(_2346_));
 sky130_fd_sc_hd__clkbuf_1 _4736_ (.A(_2346_),
    .X(_0434_));
 sky130_fd_sc_hd__a21o_1 _4737_ (.A1(\stage_gen[1].mux_gen[62].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0434_),
    .X(_0433_));
 sky130_fd_sc_hd__a21o_1 _4738_ (.A1(net29),
    .A2(_2341_),
    .B1(_0436_),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _4739_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[63].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net30),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _4740_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[63].S.IN1_L2 ),
    .X(_2347_));
 sky130_fd_sc_hd__clkbuf_1 _4741_ (.A(_2347_),
    .X(_0439_));
 sky130_fd_sc_hd__a21o_1 _4742_ (.A1(\stage_gen[1].mux_gen[63].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0439_),
    .X(_0438_));
 sky130_fd_sc_hd__a21o_1 _4743_ (.A1(net31),
    .A2(_2341_),
    .B1(_0441_),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[64].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net32),
    .X(_0442_));
 sky130_fd_sc_hd__and3_1 _4745_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[64].S.IN1_L2 ),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_1 _4746_ (.A(_2348_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _4747_ (.A1(\stage_gen[1].mux_gen[64].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0444_),
    .X(_0443_));
 sky130_fd_sc_hd__a21o_1 _4748_ (.A1(net33),
    .A2(_2341_),
    .B1(_0446_),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _4749_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[65].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net35),
    .X(_0447_));
 sky130_fd_sc_hd__and3_1 _4750_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[65].S.IN1_L2 ),
    .X(_2349_));
 sky130_fd_sc_hd__clkbuf_1 _4751_ (.A(_2349_),
    .X(_0449_));
 sky130_fd_sc_hd__a21o_1 _4752_ (.A1(\stage_gen[1].mux_gen[65].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0449_),
    .X(_0448_));
 sky130_fd_sc_hd__a21o_1 _4753_ (.A1(net36),
    .A2(_2341_),
    .B1(_0451_),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _4754_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[66].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net37),
    .X(_0452_));
 sky130_fd_sc_hd__and3_1 _4755_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[66].S.IN1_L2 ),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_1 _4756_ (.A(_2350_),
    .X(_0454_));
 sky130_fd_sc_hd__a21o_1 _4757_ (.A1(\stage_gen[1].mux_gen[66].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0454_),
    .X(_0453_));
 sky130_fd_sc_hd__a21o_1 _4758_ (.A1(net38),
    .A2(_2341_),
    .B1(_0456_),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _4759_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[67].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net39),
    .X(_0457_));
 sky130_fd_sc_hd__and3_1 _4760_ (.A(_2339_),
    .B(_2336_),
    .C(\stage_gen[1].mux_gen[67].S.IN1_L2 ),
    .X(_2351_));
 sky130_fd_sc_hd__clkbuf_1 _4761_ (.A(_2351_),
    .X(_0459_));
 sky130_fd_sc_hd__a21o_1 _4762_ (.A1(\stage_gen[1].mux_gen[67].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0459_),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_1 _4763_ (.A1(net40),
    .A2(_2341_),
    .B1(_0461_),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _4764_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[68].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net41),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_2 _4765_ (.A(_2164_),
    .X(_2352_));
 sky130_fd_sc_hd__and3_1 _4766_ (.A(_2339_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[68].S.IN1_L2 ),
    .X(_2353_));
 sky130_fd_sc_hd__clkbuf_1 _4767_ (.A(_2353_),
    .X(_0464_));
 sky130_fd_sc_hd__a21o_1 _4768_ (.A1(\stage_gen[1].mux_gen[68].S.IN1_L1 ),
    .A2(_2338_),
    .B1(_0464_),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _4769_ (.A1(net42),
    .A2(_2341_),
    .B1(_0466_),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _4770_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[69].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net43),
    .X(_0467_));
 sky130_fd_sc_hd__buf_2 _4771_ (.A(_2033_),
    .X(_2354_));
 sky130_fd_sc_hd__clkbuf_2 _4772_ (.A(_2274_),
    .X(_2355_));
 sky130_fd_sc_hd__and3_1 _4773_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[69].S.IN1_L2 ),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _4774_ (.A(_2356_),
    .X(_0469_));
 sky130_fd_sc_hd__a21o_1 _4775_ (.A1(\stage_gen[1].mux_gen[69].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0469_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_4 _4776_ (.A(_2032_),
    .X(_2357_));
 sky130_fd_sc_hd__a21o_1 _4777_ (.A1(net44),
    .A2(_2357_),
    .B1(_0471_),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _4778_ (.A1(_2343_),
    .A2(\stage_gen[1].mux_gen[70].S.IN1_L1 ),
    .B1(_2344_),
    .B2(net46),
    .X(_0477_));
 sky130_fd_sc_hd__and3_1 _4779_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[70].S.IN1_L2 ),
    .X(_2358_));
 sky130_fd_sc_hd__clkbuf_1 _4780_ (.A(_2358_),
    .X(_0479_));
 sky130_fd_sc_hd__a21o_1 _4781_ (.A1(\stage_gen[1].mux_gen[70].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0479_),
    .X(_0478_));
 sky130_fd_sc_hd__a21o_1 _4782_ (.A1(net47),
    .A2(_2357_),
    .B1(_0481_),
    .X(_0480_));
 sky130_fd_sc_hd__buf_2 _4783_ (.A(_2237_),
    .X(_2359_));
 sky130_fd_sc_hd__buf_2 _4784_ (.A(_2259_),
    .X(_2360_));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[71].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net48),
    .X(_0482_));
 sky130_fd_sc_hd__and3_1 _4786_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[71].S.IN1_L2 ),
    .X(_2361_));
 sky130_fd_sc_hd__clkbuf_1 _4787_ (.A(_2361_),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_1 _4788_ (.A1(\stage_gen[1].mux_gen[71].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0484_),
    .X(_0483_));
 sky130_fd_sc_hd__a21o_1 _4789_ (.A1(net49),
    .A2(_2357_),
    .B1(_0486_),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _4790_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[72].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net50),
    .X(_0487_));
 sky130_fd_sc_hd__and3_1 _4791_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[72].S.IN1_L2 ),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _4792_ (.A(_2362_),
    .X(_0489_));
 sky130_fd_sc_hd__a21o_1 _4793_ (.A1(\stage_gen[1].mux_gen[72].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0489_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_1 _4794_ (.A1(net51),
    .A2(_2357_),
    .B1(_0491_),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _4795_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[73].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net52),
    .X(_0492_));
 sky130_fd_sc_hd__and3_1 _4796_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[73].S.IN1_L2 ),
    .X(_2363_));
 sky130_fd_sc_hd__clkbuf_1 _4797_ (.A(_2363_),
    .X(_0494_));
 sky130_fd_sc_hd__a21o_1 _4798_ (.A1(\stage_gen[1].mux_gen[73].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0494_),
    .X(_0493_));
 sky130_fd_sc_hd__a21o_1 _4799_ (.A1(net53),
    .A2(_2357_),
    .B1(_0496_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _4800_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[74].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net54),
    .X(_0497_));
 sky130_fd_sc_hd__and3_1 _4801_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[74].S.IN1_L2 ),
    .X(_2364_));
 sky130_fd_sc_hd__clkbuf_1 _4802_ (.A(_2364_),
    .X(_0499_));
 sky130_fd_sc_hd__a21o_1 _4803_ (.A1(\stage_gen[1].mux_gen[74].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0499_),
    .X(_0498_));
 sky130_fd_sc_hd__a21o_1 _4804_ (.A1(net55),
    .A2(_2357_),
    .B1(_0501_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _4805_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[75].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net57),
    .X(_0502_));
 sky130_fd_sc_hd__and3_1 _4806_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[75].S.IN1_L2 ),
    .X(_2365_));
 sky130_fd_sc_hd__clkbuf_1 _4807_ (.A(_2365_),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_1 _4808_ (.A1(\stage_gen[1].mux_gen[75].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0504_),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _4809_ (.A1(net58),
    .A2(_2357_),
    .B1(_0506_),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _4810_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[76].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net59),
    .X(_0507_));
 sky130_fd_sc_hd__and3_1 _4811_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[76].S.IN1_L2 ),
    .X(_2366_));
 sky130_fd_sc_hd__clkbuf_1 _4812_ (.A(_2366_),
    .X(_0509_));
 sky130_fd_sc_hd__a21o_1 _4813_ (.A1(\stage_gen[1].mux_gen[76].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0509_),
    .X(_0508_));
 sky130_fd_sc_hd__a21o_1 _4814_ (.A1(net60),
    .A2(_2357_),
    .B1(_0511_),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _4815_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[77].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net61),
    .X(_0512_));
 sky130_fd_sc_hd__and3_1 _4816_ (.A(_2355_),
    .B(_2352_),
    .C(\stage_gen[1].mux_gen[77].S.IN1_L2 ),
    .X(_2367_));
 sky130_fd_sc_hd__clkbuf_1 _4817_ (.A(_2367_),
    .X(_0514_));
 sky130_fd_sc_hd__a21o_1 _4818_ (.A1(\stage_gen[1].mux_gen[77].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0514_),
    .X(_0513_));
 sky130_fd_sc_hd__a21o_1 _4819_ (.A1(net62),
    .A2(_2357_),
    .B1(_0516_),
    .X(_0515_));
 sky130_fd_sc_hd__a22o_1 _4820_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[78].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net63),
    .X(_0517_));
 sky130_fd_sc_hd__buf_2 _4821_ (.A(_1377_),
    .X(_2368_));
 sky130_fd_sc_hd__and3_1 _4822_ (.A(_2355_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[78].S.IN1_L2 ),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _4823_ (.A(_2369_),
    .X(_0519_));
 sky130_fd_sc_hd__a21o_1 _4824_ (.A1(\stage_gen[1].mux_gen[78].S.IN1_L1 ),
    .A2(_2354_),
    .B1(_0519_),
    .X(_0518_));
 sky130_fd_sc_hd__a21o_1 _4825_ (.A1(net64),
    .A2(_2357_),
    .B1(_0521_),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _4826_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[79].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net65),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _4827_ (.A(_2033_),
    .X(_2370_));
 sky130_fd_sc_hd__clkbuf_2 _4828_ (.A(_2274_),
    .X(_2371_));
 sky130_fd_sc_hd__and3_1 _4829_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[79].S.IN1_L2 ),
    .X(_2372_));
 sky130_fd_sc_hd__buf_6 _4830_ (.A(_2372_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _4831_ (.A1(\stage_gen[1].mux_gen[79].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0524_),
    .X(_0523_));
 sky130_fd_sc_hd__buf_4 _4832_ (.A(_2032_),
    .X(_2373_));
 sky130_fd_sc_hd__a21o_1 _4833_ (.A1(net66),
    .A2(_2373_),
    .B1(_0526_),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _4834_ (.A1(_2359_),
    .A2(\stage_gen[1].mux_gen[80].S.IN1_L1 ),
    .B1(_2360_),
    .B2(net68),
    .X(_0532_));
 sky130_fd_sc_hd__and3_1 _4835_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[80].S.IN1_L2 ),
    .X(_2374_));
 sky130_fd_sc_hd__clkbuf_1 _4836_ (.A(_2374_),
    .X(_0534_));
 sky130_fd_sc_hd__a21o_1 _4837_ (.A1(\stage_gen[1].mux_gen[80].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0534_),
    .X(_0533_));
 sky130_fd_sc_hd__a21o_1 _4838_ (.A1(net69),
    .A2(_2373_),
    .B1(_0536_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_4 _4839_ (.A(_2237_),
    .X(_2375_));
 sky130_fd_sc_hd__clkbuf_4 _4840_ (.A(_2259_),
    .X(_2376_));
 sky130_fd_sc_hd__a22o_1 _4841_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[81].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net70),
    .X(_0537_));
 sky130_fd_sc_hd__and3_1 _4842_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[81].S.IN1_L2 ),
    .X(_2377_));
 sky130_fd_sc_hd__clkbuf_1 _4843_ (.A(_2377_),
    .X(_0539_));
 sky130_fd_sc_hd__a21o_1 _4844_ (.A1(\stage_gen[1].mux_gen[81].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0539_),
    .X(_0538_));
 sky130_fd_sc_hd__a21o_1 _4845_ (.A1(net71),
    .A2(_2373_),
    .B1(_0541_),
    .X(_0540_));
 sky130_fd_sc_hd__a22o_1 _4846_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[82].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net72),
    .X(_0542_));
 sky130_fd_sc_hd__and3_1 _4847_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[82].S.IN1_L2 ),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _4848_ (.A(_2378_),
    .X(_0544_));
 sky130_fd_sc_hd__a21o_1 _4849_ (.A1(\stage_gen[1].mux_gen[82].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0544_),
    .X(_0543_));
 sky130_fd_sc_hd__a21o_1 _4850_ (.A1(net73),
    .A2(_2373_),
    .B1(_0546_),
    .X(_0545_));
 sky130_fd_sc_hd__a22o_1 _4851_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[83].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net74),
    .X(_0547_));
 sky130_fd_sc_hd__and3_1 _4852_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[83].S.IN1_L2 ),
    .X(_2379_));
 sky130_fd_sc_hd__clkbuf_1 _4853_ (.A(_2379_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _4854_ (.A1(\stage_gen[1].mux_gen[83].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0549_),
    .X(_0548_));
 sky130_fd_sc_hd__a21o_1 _4855_ (.A1(net75),
    .A2(_2373_),
    .B1(_0551_),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _4856_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[84].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net76),
    .X(_0552_));
 sky130_fd_sc_hd__and3_1 _4857_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[84].S.IN1_L2 ),
    .X(_2380_));
 sky130_fd_sc_hd__clkbuf_1 _4858_ (.A(_2380_),
    .X(_0554_));
 sky130_fd_sc_hd__a21o_1 _4859_ (.A1(\stage_gen[1].mux_gen[84].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0554_),
    .X(_0553_));
 sky130_fd_sc_hd__a21o_1 _4860_ (.A1(net77),
    .A2(_2373_),
    .B1(_0556_),
    .X(_0555_));
 sky130_fd_sc_hd__a22o_1 _4861_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[85].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net79),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _4862_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[85].S.IN1_L2 ),
    .X(_2381_));
 sky130_fd_sc_hd__clkbuf_1 _4863_ (.A(_2381_),
    .X(_0559_));
 sky130_fd_sc_hd__a21o_1 _4864_ (.A1(\stage_gen[1].mux_gen[85].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0559_),
    .X(_0558_));
 sky130_fd_sc_hd__a21o_1 _4865_ (.A1(net80),
    .A2(_2373_),
    .B1(_0561_),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _4866_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[86].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net81),
    .X(_0562_));
 sky130_fd_sc_hd__and3_1 _4867_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[86].S.IN1_L2 ),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _4868_ (.A(_2382_),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _4869_ (.A1(\stage_gen[1].mux_gen[86].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0564_),
    .X(_0563_));
 sky130_fd_sc_hd__a21o_1 _4870_ (.A1(net82),
    .A2(_2373_),
    .B1(_0566_),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _4871_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[87].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net83),
    .X(_0567_));
 sky130_fd_sc_hd__and3_1 _4872_ (.A(_2371_),
    .B(_2368_),
    .C(\stage_gen[1].mux_gen[87].S.IN1_L2 ),
    .X(_2383_));
 sky130_fd_sc_hd__clkbuf_1 _4873_ (.A(_2383_),
    .X(_0569_));
 sky130_fd_sc_hd__a21o_1 _4874_ (.A1(\stage_gen[1].mux_gen[87].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0569_),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_1 _4875_ (.A1(net84),
    .A2(_2373_),
    .B1(_0571_),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _4876_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[88].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net85),
    .X(_0572_));
 sky130_fd_sc_hd__buf_2 _4877_ (.A(_1377_),
    .X(_2384_));
 sky130_fd_sc_hd__and3_1 _4878_ (.A(_2371_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[88].S.IN1_L2 ),
    .X(_2385_));
 sky130_fd_sc_hd__clkbuf_1 _4879_ (.A(_2385_),
    .X(_0574_));
 sky130_fd_sc_hd__a21o_1 _4880_ (.A1(\stage_gen[1].mux_gen[88].S.IN1_L1 ),
    .A2(_2370_),
    .B1(_0574_),
    .X(_0573_));
 sky130_fd_sc_hd__a21o_1 _4881_ (.A1(net86),
    .A2(_2373_),
    .B1(_0576_),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _4882_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[89].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net87),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_4 _4883_ (.A(_2033_),
    .X(_2386_));
 sky130_fd_sc_hd__clkbuf_2 _4884_ (.A(_2274_),
    .X(_2387_));
 sky130_fd_sc_hd__and3_1 _4885_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[89].S.IN1_L2 ),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _4886_ (.A(_2388_),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_1 _4887_ (.A1(\stage_gen[1].mux_gen[89].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0579_),
    .X(_0578_));
 sky130_fd_sc_hd__buf_4 _4888_ (.A(_2032_),
    .X(_2389_));
 sky130_fd_sc_hd__a21o_1 _4889_ (.A1(net88),
    .A2(_2389_),
    .B1(_0581_),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _4890_ (.A1(_2375_),
    .A2(\stage_gen[1].mux_gen[90].S.IN1_L1 ),
    .B1(_2376_),
    .B2(net90),
    .X(_0587_));
 sky130_fd_sc_hd__and3_1 _4891_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[90].S.IN1_L2 ),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _4892_ (.A(_2390_),
    .X(_0589_));
 sky130_fd_sc_hd__a21o_1 _4893_ (.A1(\stage_gen[1].mux_gen[90].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0589_),
    .X(_0588_));
 sky130_fd_sc_hd__a21o_1 _4894_ (.A1(net91),
    .A2(_2389_),
    .B1(_0591_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_4 _4895_ (.A(_2237_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_4 _4896_ (.A(_2259_),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _4897_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[91].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net92),
    .X(_0592_));
 sky130_fd_sc_hd__and3_1 _4898_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[91].S.IN1_L2 ),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _4899_ (.A(_2393_),
    .X(_0594_));
 sky130_fd_sc_hd__a21o_1 _4900_ (.A1(\stage_gen[1].mux_gen[91].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0594_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _4901_ (.A1(net93),
    .A2(_2389_),
    .B1(_0596_),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _4902_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[92].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net94),
    .X(_0597_));
 sky130_fd_sc_hd__and3_1 _4903_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[92].S.IN1_L2 ),
    .X(_2394_));
 sky130_fd_sc_hd__clkbuf_1 _4904_ (.A(_2394_),
    .X(_0599_));
 sky130_fd_sc_hd__a21o_1 _4905_ (.A1(\stage_gen[1].mux_gen[92].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0599_),
    .X(_0598_));
 sky130_fd_sc_hd__a21o_1 _4906_ (.A1(net95),
    .A2(_2389_),
    .B1(_0601_),
    .X(_0600_));
 sky130_fd_sc_hd__a22o_1 _4907_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[93].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net96),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _4908_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[93].S.IN1_L2 ),
    .X(_2395_));
 sky130_fd_sc_hd__clkbuf_1 _4909_ (.A(_2395_),
    .X(_0604_));
 sky130_fd_sc_hd__a21o_1 _4910_ (.A1(\stage_gen[1].mux_gen[93].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0604_),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _4911_ (.A1(net97),
    .A2(_2389_),
    .B1(_0606_),
    .X(_0605_));
 sky130_fd_sc_hd__a22o_1 _4912_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[94].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net98),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _4913_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[94].S.IN1_L2 ),
    .X(_2396_));
 sky130_fd_sc_hd__clkbuf_1 _4914_ (.A(_2396_),
    .X(_0609_));
 sky130_fd_sc_hd__a21o_1 _4915_ (.A1(\stage_gen[1].mux_gen[94].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0609_),
    .X(_0608_));
 sky130_fd_sc_hd__a21o_1 _4916_ (.A1(net99),
    .A2(_2389_),
    .B1(_0611_),
    .X(_0610_));
 sky130_fd_sc_hd__a22o_1 _4917_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[95].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net101),
    .X(_0612_));
 sky130_fd_sc_hd__and3_1 _4918_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[95].S.IN1_L2 ),
    .X(_2397_));
 sky130_fd_sc_hd__clkbuf_1 _4919_ (.A(_2397_),
    .X(_0614_));
 sky130_fd_sc_hd__a21o_1 _4920_ (.A1(\stage_gen[1].mux_gen[95].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0614_),
    .X(_0613_));
 sky130_fd_sc_hd__a21o_1 _4921_ (.A1(net102),
    .A2(_2389_),
    .B1(_0616_),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_1 _4922_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[96].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net103),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _4923_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[96].S.IN1_L2 ),
    .X(_2398_));
 sky130_fd_sc_hd__buf_6 _4924_ (.A(_2398_),
    .X(_0619_));
 sky130_fd_sc_hd__a21o_1 _4925_ (.A1(\stage_gen[1].mux_gen[96].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0619_),
    .X(_0618_));
 sky130_fd_sc_hd__a21o_1 _4926_ (.A1(net104),
    .A2(_2389_),
    .B1(_0621_),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _4927_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[97].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net105),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _4928_ (.A(_2387_),
    .B(_2384_),
    .C(\stage_gen[1].mux_gen[97].S.IN1_L2 ),
    .X(_2399_));
 sky130_fd_sc_hd__clkbuf_1 _4929_ (.A(_2399_),
    .X(_0624_));
 sky130_fd_sc_hd__a21o_1 _4930_ (.A1(\stage_gen[1].mux_gen[97].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0624_),
    .X(_0623_));
 sky130_fd_sc_hd__a21o_1 _4931_ (.A1(net106),
    .A2(_2389_),
    .B1(_0626_),
    .X(_0625_));
 sky130_fd_sc_hd__a22o_1 _4932_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[98].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net107),
    .X(_0627_));
 sky130_fd_sc_hd__buf_2 _4933_ (.A(_1377_),
    .X(_2400_));
 sky130_fd_sc_hd__and3_1 _4934_ (.A(_2387_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[98].S.IN1_L2 ),
    .X(_2401_));
 sky130_fd_sc_hd__clkbuf_1 _4935_ (.A(_2401_),
    .X(_0629_));
 sky130_fd_sc_hd__a21o_1 _4936_ (.A1(\stage_gen[1].mux_gen[98].S.IN1_L1 ),
    .A2(_2386_),
    .B1(_0629_),
    .X(_0628_));
 sky130_fd_sc_hd__a21o_1 _4937_ (.A1(net108),
    .A2(_2389_),
    .B1(_0631_),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _4938_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[99].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net109),
    .X(_0632_));
 sky130_fd_sc_hd__buf_4 _4939_ (.A(_2033_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_4 _4940_ (.A(_2274_),
    .X(_2403_));
 sky130_fd_sc_hd__and3_1 _4941_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[99].S.IN1_L2 ),
    .X(_2404_));
 sky130_fd_sc_hd__clkbuf_1 _4942_ (.A(_2404_),
    .X(_0634_));
 sky130_fd_sc_hd__a21o_1 _4943_ (.A1(\stage_gen[1].mux_gen[99].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0634_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _4944_ (.A(_2032_),
    .X(_2405_));
 sky130_fd_sc_hd__a21o_1 _4945_ (.A1(net110),
    .A2(_2405_),
    .B1(_0636_),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_1 _4946_ (.A1(_2391_),
    .A2(\stage_gen[1].mux_gen[100].S.IN1_L1 ),
    .B1(_2392_),
    .B2(net113),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _4947_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[100].S.IN1_L2 ),
    .X(_2406_));
 sky130_fd_sc_hd__clkbuf_1 _4948_ (.A(_2406_),
    .X(_0009_));
 sky130_fd_sc_hd__a21o_1 _4949_ (.A1(\stage_gen[1].mux_gen[100].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0009_),
    .X(_0008_));
 sky130_fd_sc_hd__a21o_1 _4950_ (.A1(net114),
    .A2(_2405_),
    .B1(_0011_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_4 _4951_ (.A(_2237_),
    .X(_2407_));
 sky130_fd_sc_hd__buf_4 _4952_ (.A(_2259_),
    .X(_2408_));
 sky130_fd_sc_hd__a22o_1 _4953_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[101].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net115),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _4954_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[101].S.IN1_L2 ),
    .X(_2409_));
 sky130_fd_sc_hd__clkbuf_1 _4955_ (.A(_2409_),
    .X(_0014_));
 sky130_fd_sc_hd__a21o_1 _4956_ (.A1(\stage_gen[1].mux_gen[101].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0014_),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _4957_ (.A1(net116),
    .A2(_2405_),
    .B1(_0016_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _4958_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[102].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net117),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _4959_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[102].S.IN1_L2 ),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_1 _4960_ (.A(_2410_),
    .X(_0019_));
 sky130_fd_sc_hd__a21o_1 _4961_ (.A1(\stage_gen[1].mux_gen[102].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0019_),
    .X(_0018_));
 sky130_fd_sc_hd__a21o_1 _4962_ (.A1(net118),
    .A2(_2405_),
    .B1(_0021_),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _4963_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[103].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net119),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _4964_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[103].S.IN1_L2 ),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _4965_ (.A(_2411_),
    .X(_0024_));
 sky130_fd_sc_hd__a21o_1 _4966_ (.A1(\stage_gen[1].mux_gen[103].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0024_),
    .X(_0023_));
 sky130_fd_sc_hd__a21o_1 _4967_ (.A1(net120),
    .A2(_2405_),
    .B1(_0026_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _4968_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[104].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net121),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _4969_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[104].S.IN1_L2 ),
    .X(_2412_));
 sky130_fd_sc_hd__clkbuf_1 _4970_ (.A(_2412_),
    .X(_0029_));
 sky130_fd_sc_hd__a21o_1 _4971_ (.A1(\stage_gen[1].mux_gen[104].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0029_),
    .X(_0028_));
 sky130_fd_sc_hd__a21o_1 _4972_ (.A1(net122),
    .A2(_2405_),
    .B1(_0031_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _4973_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[105].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net124),
    .X(_0032_));
 sky130_fd_sc_hd__and3_1 _4974_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[105].S.IN1_L2 ),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _4975_ (.A(_2413_),
    .X(_0034_));
 sky130_fd_sc_hd__a21o_1 _4976_ (.A1(\stage_gen[1].mux_gen[105].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0034_),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _4977_ (.A1(net125),
    .A2(_2405_),
    .B1(_0036_),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _4978_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[106].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net126),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _4979_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[106].S.IN1_L2 ),
    .X(_2414_));
 sky130_fd_sc_hd__clkbuf_1 _4980_ (.A(_2414_),
    .X(_0039_));
 sky130_fd_sc_hd__a21o_1 _4981_ (.A1(\stage_gen[1].mux_gen[106].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0039_),
    .X(_0038_));
 sky130_fd_sc_hd__a21o_1 _4982_ (.A1(net127),
    .A2(_2405_),
    .B1(_0041_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _4983_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[107].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net128),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _4984_ (.A(_2403_),
    .B(_2400_),
    .C(\stage_gen[1].mux_gen[107].S.IN1_L2 ),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_1 _4985_ (.A(_2415_),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _4986_ (.A1(\stage_gen[1].mux_gen[107].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0044_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _4987_ (.A1(net129),
    .A2(_2405_),
    .B1(_0046_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _4988_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[108].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net130),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _4989_ (.A(_1377_),
    .X(_2416_));
 sky130_fd_sc_hd__and3_1 _4990_ (.A(_2403_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[108].S.IN1_L2 ),
    .X(_2417_));
 sky130_fd_sc_hd__clkbuf_1 _4991_ (.A(_2417_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _4992_ (.A1(\stage_gen[1].mux_gen[108].S.IN1_L1 ),
    .A2(_2402_),
    .B1(_0049_),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _4993_ (.A1(net131),
    .A2(_2405_),
    .B1(_0051_),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _4994_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[109].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net132),
    .X(_0052_));
 sky130_fd_sc_hd__buf_4 _4995_ (.A(_2033_),
    .X(_2418_));
 sky130_fd_sc_hd__buf_2 _4996_ (.A(_2274_),
    .X(_2419_));
 sky130_fd_sc_hd__and3_1 _4997_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[109].S.IN1_L2 ),
    .X(_2420_));
 sky130_fd_sc_hd__clkbuf_1 _4998_ (.A(_2420_),
    .X(_0054_));
 sky130_fd_sc_hd__a21o_1 _4999_ (.A1(\stage_gen[1].mux_gen[109].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0054_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_4 _5000_ (.A(_2032_),
    .X(_2421_));
 sky130_fd_sc_hd__a21o_1 _5001_ (.A1(net133),
    .A2(_2421_),
    .B1(_0056_),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _5002_ (.A1(_2407_),
    .A2(\stage_gen[1].mux_gen[110].S.IN1_L1 ),
    .B1(_2408_),
    .B2(net135),
    .X(_0062_));
 sky130_fd_sc_hd__and3_1 _5003_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[110].S.IN1_L2 ),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _5004_ (.A(_2422_),
    .X(_0064_));
 sky130_fd_sc_hd__a21o_1 _5005_ (.A1(\stage_gen[1].mux_gen[110].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0064_),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_1 _5006_ (.A1(net136),
    .A2(_2421_),
    .B1(_0066_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_4 _5007_ (.A(_2237_),
    .X(_2423_));
 sky130_fd_sc_hd__buf_4 _5008_ (.A(_2259_),
    .X(_2424_));
 sky130_fd_sc_hd__a22o_1 _5009_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[111].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net137),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _5010_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[111].S.IN1_L2 ),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _5011_ (.A(_2425_),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _5012_ (.A1(\stage_gen[1].mux_gen[111].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0069_),
    .X(_0068_));
 sky130_fd_sc_hd__a21o_1 _5013_ (.A1(net138),
    .A2(_2421_),
    .B1(_0071_),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _5014_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[112].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net139),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _5015_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[112].S.IN1_L2 ),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5016_ (.A(_2426_),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _5017_ (.A1(\stage_gen[1].mux_gen[112].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0074_),
    .X(_0073_));
 sky130_fd_sc_hd__a21o_1 _5018_ (.A1(net140),
    .A2(_2421_),
    .B1(_0076_),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _5019_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[113].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net141),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _5020_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[113].S.IN1_L2 ),
    .X(_2427_));
 sky130_fd_sc_hd__clkbuf_1 _5021_ (.A(_2427_),
    .X(_0079_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(\stage_gen[1].mux_gen[113].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0079_),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_1 _5023_ (.A1(net142),
    .A2(_2421_),
    .B1(_0081_),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _5024_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[114].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net143),
    .X(_0082_));
 sky130_fd_sc_hd__and3_1 _5025_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[114].S.IN1_L2 ),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _5026_ (.A(_2428_),
    .X(_0084_));
 sky130_fd_sc_hd__a21o_1 _5027_ (.A1(\stage_gen[1].mux_gen[114].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0084_),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _5028_ (.A1(net144),
    .A2(_2421_),
    .B1(_0086_),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _5029_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[115].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net146),
    .X(_0087_));
 sky130_fd_sc_hd__and3_1 _5030_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[115].S.IN1_L2 ),
    .X(_2429_));
 sky130_fd_sc_hd__clkbuf_1 _5031_ (.A(_2429_),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_1 _5032_ (.A1(\stage_gen[1].mux_gen[115].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0089_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _5033_ (.A1(net147),
    .A2(_2421_),
    .B1(_0091_),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _5034_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[116].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net148),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _5035_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[116].S.IN1_L2 ),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _5036_ (.A(_2430_),
    .X(_0094_));
 sky130_fd_sc_hd__a21o_1 _5037_ (.A1(\stage_gen[1].mux_gen[116].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0094_),
    .X(_0093_));
 sky130_fd_sc_hd__a21o_1 _5038_ (.A1(net149),
    .A2(_2421_),
    .B1(_0096_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _5039_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[117].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net150),
    .X(_0097_));
 sky130_fd_sc_hd__and3_1 _5040_ (.A(_2419_),
    .B(_2416_),
    .C(\stage_gen[1].mux_gen[117].S.IN1_L2 ),
    .X(_2431_));
 sky130_fd_sc_hd__clkbuf_1 _5041_ (.A(_2431_),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_1 _5042_ (.A1(\stage_gen[1].mux_gen[117].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0099_),
    .X(_0098_));
 sky130_fd_sc_hd__a21o_1 _5043_ (.A1(net151),
    .A2(_2421_),
    .B1(_0101_),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _5044_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[118].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net152),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _5045_ (.A(_1377_),
    .X(_2432_));
 sky130_fd_sc_hd__and3_1 _5046_ (.A(_2419_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[118].S.IN1_L2 ),
    .X(_2433_));
 sky130_fd_sc_hd__clkbuf_1 _5047_ (.A(_2433_),
    .X(_0104_));
 sky130_fd_sc_hd__a21o_1 _5048_ (.A1(\stage_gen[1].mux_gen[118].S.IN1_L1 ),
    .A2(_2418_),
    .B1(_0104_),
    .X(_0103_));
 sky130_fd_sc_hd__a21o_1 _5049_ (.A1(net153),
    .A2(_2421_),
    .B1(_0106_),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _5050_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[119].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net154),
    .X(_0107_));
 sky130_fd_sc_hd__and3_1 _5051_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[119].S.IN1_L2 ),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _5052_ (.A(_2434_),
    .X(_0109_));
 sky130_fd_sc_hd__a21o_1 _5053_ (.A1(\stage_gen[1].mux_gen[119].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0109_),
    .X(_0108_));
 sky130_fd_sc_hd__a21o_1 _5054_ (.A1(net155),
    .A2(_2239_),
    .B1(_0111_),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _5055_ (.A1(_2423_),
    .A2(\stage_gen[1].mux_gen[120].S.IN1_L1 ),
    .B1(_2424_),
    .B2(net157),
    .X(_0117_));
 sky130_fd_sc_hd__and3_1 _5056_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[120].S.IN1_L2 ),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _5057_ (.A(_2435_),
    .X(_0119_));
 sky130_fd_sc_hd__a21o_1 _5058_ (.A1(\stage_gen[1].mux_gen[120].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0119_),
    .X(_0118_));
 sky130_fd_sc_hd__a21o_1 _5059_ (.A1(net158),
    .A2(_2239_),
    .B1(_0121_),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _5060_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[121].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net159),
    .X(_0122_));
 sky130_fd_sc_hd__and3_1 _5061_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[121].S.IN1_L2 ),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5062_ (.A(_2436_),
    .X(_0124_));
 sky130_fd_sc_hd__a21o_1 _5063_ (.A1(\stage_gen[1].mux_gen[121].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0124_),
    .X(_0123_));
 sky130_fd_sc_hd__a21o_1 _5064_ (.A1(net160),
    .A2(_2239_),
    .B1(_0126_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _5065_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[122].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net161),
    .X(_0127_));
 sky130_fd_sc_hd__and3_1 _5066_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[122].S.IN1_L2 ),
    .X(_2437_));
 sky130_fd_sc_hd__clkbuf_1 _5067_ (.A(_2437_),
    .X(_0129_));
 sky130_fd_sc_hd__a21o_1 _5068_ (.A1(\stage_gen[1].mux_gen[122].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0129_),
    .X(_0128_));
 sky130_fd_sc_hd__a21o_1 _5069_ (.A1(net162),
    .A2(_2239_),
    .B1(_0131_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _5070_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[123].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net163),
    .X(_0132_));
 sky130_fd_sc_hd__and3_1 _5071_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[123].S.IN1_L2 ),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_1 _5072_ (.A(_2438_),
    .X(_0134_));
 sky130_fd_sc_hd__a21o_1 _5073_ (.A1(\stage_gen[1].mux_gen[123].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0134_),
    .X(_0133_));
 sky130_fd_sc_hd__a21o_1 _5074_ (.A1(net164),
    .A2(_2239_),
    .B1(_0136_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _5075_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[124].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net165),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _5076_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[124].S.IN1_L2 ),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _5077_ (.A(_2439_),
    .X(_0139_));
 sky130_fd_sc_hd__a21o_1 _5078_ (.A1(\stage_gen[1].mux_gen[124].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0139_),
    .X(_0138_));
 sky130_fd_sc_hd__a21o_1 _5079_ (.A1(net166),
    .A2(_2239_),
    .B1(_0141_),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _5080_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[125].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net168),
    .X(_0142_));
 sky130_fd_sc_hd__and3_1 _5081_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[125].S.IN1_L2 ),
    .X(_2440_));
 sky130_fd_sc_hd__clkbuf_1 _5082_ (.A(_2440_),
    .X(_0144_));
 sky130_fd_sc_hd__a21o_1 _5083_ (.A1(\stage_gen[1].mux_gen[125].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0144_),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _5084_ (.A1(net169),
    .A2(_2239_),
    .B1(_0146_),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _5085_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[126].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net170),
    .X(_0147_));
 sky130_fd_sc_hd__and3_1 _5086_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[126].S.IN1_L2 ),
    .X(_2441_));
 sky130_fd_sc_hd__clkbuf_1 _5087_ (.A(_2441_),
    .X(_0149_));
 sky130_fd_sc_hd__a21o_1 _5088_ (.A1(\stage_gen[1].mux_gen[126].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0149_),
    .X(_0148_));
 sky130_fd_sc_hd__a21o_1 _5089_ (.A1(net171),
    .A2(_2239_),
    .B1(_0151_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _5090_ (.A1(_1370_),
    .A2(\stage_gen[1].mux_gen[127].S.IN1_L1 ),
    .B1(_1375_),
    .B2(net172),
    .X(_0152_));
 sky130_fd_sc_hd__and3_1 _5091_ (.A(_2256_),
    .B(_2432_),
    .C(\stage_gen[1].mux_gen[127].S.IN1_L2 ),
    .X(_2442_));
 sky130_fd_sc_hd__clkbuf_1 _5092_ (.A(_2442_),
    .X(_0154_));
 sky130_fd_sc_hd__a21o_1 _5093_ (.A1(\stage_gen[1].mux_gen[127].S.IN1_L1 ),
    .A2(_2238_),
    .B1(_0154_),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_1 _5094_ (.A1(net173),
    .A2(_2239_),
    .B1(_0156_),
    .X(_0155_));
 sky130_fd_sc_hd__buf_4 _5095_ (.A(_1421_),
    .X(_2443_));
 sky130_fd_sc_hd__a22oi_1 _5096_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[0].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[0].S.IN1_L3 ),
    .Y(_2444_));
 sky130_fd_sc_hd__clkbuf_4 _5097_ (.A(_1387_),
    .X(_2445_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[0].S.IN1_L1 ),
    .Y(_2446_));
 sky130_fd_sc_hd__o21ai_1 _5099_ (.A1(_2443_),
    .A2(_2444_),
    .B1(_2446_),
    .Y(_0642_));
 sky130_fd_sc_hd__and3_1 _5100_ (.A(_1517_),
    .B(_1961_),
    .C(\stage_gen[2].mux_gen[0].S.IN1_L2 ),
    .X(_2447_));
 sky130_fd_sc_hd__clkbuf_1 _5101_ (.A(_2447_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2b_1 _5102_ (.A_N(_0644_),
    .B(_2446_),
    .Y(_2448_));
 sky130_fd_sc_hd__clkbuf_1 _5103_ (.A(_2448_),
    .X(_0643_));
 sky130_fd_sc_hd__a22oi_1 _5104_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[1].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[1].S.IN1_L3 ),
    .Y(_2449_));
 sky130_fd_sc_hd__o21bai_1 _5105_ (.A1(_1529_),
    .A2(_2449_),
    .B1_N(_0646_),
    .Y(_0645_));
 sky130_fd_sc_hd__a22oi_1 _5106_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[2].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[2].S.IN1_L3 ),
    .Y(_2450_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[1].S.IN1_L1 ),
    .Y(_2451_));
 sky130_fd_sc_hd__o21ai_1 _5108_ (.A1(_2443_),
    .A2(_2450_),
    .B1(_2451_),
    .Y(_0699_));
 sky130_fd_sc_hd__clkbuf_4 _5109_ (.A(_1384_),
    .X(_2452_));
 sky130_fd_sc_hd__and3_1 _5110_ (.A(_1517_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[1].S.IN1_L2 ),
    .X(_2453_));
 sky130_fd_sc_hd__clkbuf_1 _5111_ (.A(_2453_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2b_1 _5112_ (.A_N(_0701_),
    .B(_2451_),
    .Y(_2454_));
 sky130_fd_sc_hd__clkbuf_1 _5113_ (.A(_2454_),
    .X(_0700_));
 sky130_fd_sc_hd__a22oi_1 _5114_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[3].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[3].S.IN1_L3 ),
    .Y(_2455_));
 sky130_fd_sc_hd__o21bai_1 _5115_ (.A1(_1529_),
    .A2(_2455_),
    .B1_N(_0703_),
    .Y(_0702_));
 sky130_fd_sc_hd__a22oi_1 _5116_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[4].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[4].S.IN1_L3 ),
    .Y(_2456_));
 sky130_fd_sc_hd__nand2_1 _5117_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[2].S.IN1_L1 ),
    .Y(_2457_));
 sky130_fd_sc_hd__o21ai_1 _5118_ (.A1(_2443_),
    .A2(_2456_),
    .B1(_2457_),
    .Y(_0754_));
 sky130_fd_sc_hd__and3_1 _5119_ (.A(_1517_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[2].S.IN1_L2 ),
    .X(_2458_));
 sky130_fd_sc_hd__clkbuf_1 _5120_ (.A(_2458_),
    .X(_0756_));
 sky130_fd_sc_hd__nand2b_1 _5121_ (.A_N(_0756_),
    .B(_2457_),
    .Y(_2459_));
 sky130_fd_sc_hd__clkbuf_1 _5122_ (.A(_2459_),
    .X(_0755_));
 sky130_fd_sc_hd__a22oi_1 _5123_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[5].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[5].S.IN1_L3 ),
    .Y(_2460_));
 sky130_fd_sc_hd__o21bai_1 _5124_ (.A1(_1529_),
    .A2(_2460_),
    .B1_N(_0758_),
    .Y(_0757_));
 sky130_fd_sc_hd__a22oi_1 _5125_ (.A1(_1522_),
    .A2(\stage_gen[1].mux_gen[6].S.IN1_L5 ),
    .B1(_1523_),
    .B2(\stage_gen[1].mux_gen[6].S.IN1_L3 ),
    .Y(_2461_));
 sky130_fd_sc_hd__nand2_1 _5126_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[3].S.IN1_L1 ),
    .Y(_2462_));
 sky130_fd_sc_hd__o21ai_1 _5127_ (.A1(_2443_),
    .A2(_2461_),
    .B1(_2462_),
    .Y(_0809_));
 sky130_fd_sc_hd__buf_2 _5128_ (.A(_1445_),
    .X(_2463_));
 sky130_fd_sc_hd__and3_1 _5129_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[3].S.IN1_L2 ),
    .X(_2464_));
 sky130_fd_sc_hd__clkbuf_1 _5130_ (.A(_2464_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2b_1 _5131_ (.A_N(_0811_),
    .B(_2462_),
    .Y(_2465_));
 sky130_fd_sc_hd__clkbuf_1 _5132_ (.A(_2465_),
    .X(_0810_));
 sky130_fd_sc_hd__a22oi_1 _5133_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[7].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[7].S.IN1_L3 ),
    .Y(_2466_));
 sky130_fd_sc_hd__o21bai_1 _5134_ (.A1(_1529_),
    .A2(_2466_),
    .B1_N(_0813_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_4 _5135_ (.A(_1368_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_4 _5136_ (.A(_1373_),
    .X(_2468_));
 sky130_fd_sc_hd__a22oi_1 _5137_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[8].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[8].S.IN1_L3 ),
    .Y(_2469_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[4].S.IN1_L1 ),
    .Y(_2470_));
 sky130_fd_sc_hd__o21ai_1 _5139_ (.A1(_2443_),
    .A2(_2469_),
    .B1(_2470_),
    .Y(_0864_));
 sky130_fd_sc_hd__and3_1 _5140_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[4].S.IN1_L2 ),
    .X(_2471_));
 sky130_fd_sc_hd__clkbuf_1 _5141_ (.A(_2471_),
    .X(_0866_));
 sky130_fd_sc_hd__nand2b_1 _5142_ (.A_N(_0866_),
    .B(_2470_),
    .Y(_2472_));
 sky130_fd_sc_hd__clkbuf_1 _5143_ (.A(_2472_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_4 _5144_ (.A(_1421_),
    .X(_2473_));
 sky130_fd_sc_hd__a22oi_1 _5145_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[9].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[9].S.IN1_L3 ),
    .Y(_2474_));
 sky130_fd_sc_hd__o21bai_1 _5146_ (.A1(_2473_),
    .A2(_2474_),
    .B1_N(_0868_),
    .Y(_0867_));
 sky130_fd_sc_hd__a22oi_2 _5147_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[10].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[10].S.IN1_L3 ),
    .Y(_2475_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[5].S.IN1_L1 ),
    .Y(_2476_));
 sky130_fd_sc_hd__o21ai_1 _5149_ (.A1(_2443_),
    .A2(_2475_),
    .B1(_2476_),
    .Y(_0919_));
 sky130_fd_sc_hd__and3_1 _5150_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[5].S.IN1_L2 ),
    .X(_2477_));
 sky130_fd_sc_hd__clkbuf_1 _5151_ (.A(_2477_),
    .X(_0921_));
 sky130_fd_sc_hd__nand2b_1 _5152_ (.A_N(_0921_),
    .B(_2476_),
    .Y(_2478_));
 sky130_fd_sc_hd__clkbuf_1 _5153_ (.A(_2478_),
    .X(_0920_));
 sky130_fd_sc_hd__a22oi_1 _5154_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[11].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[11].S.IN1_L3 ),
    .Y(_2479_));
 sky130_fd_sc_hd__o21bai_1 _5155_ (.A1(_2473_),
    .A2(_2479_),
    .B1_N(_0923_),
    .Y(_0922_));
 sky130_fd_sc_hd__a22oi_1 _5156_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[12].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[12].S.IN1_L3 ),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[6].S.IN1_L1 ),
    .Y(_2481_));
 sky130_fd_sc_hd__o21ai_1 _5158_ (.A1(_2443_),
    .A2(_2480_),
    .B1(_2481_),
    .Y(_0944_));
 sky130_fd_sc_hd__and3_1 _5159_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[6].S.IN1_L2 ),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _5160_ (.A(_2482_),
    .X(_0946_));
 sky130_fd_sc_hd__nand2b_1 _5161_ (.A_N(_0946_),
    .B(_2481_),
    .Y(_2483_));
 sky130_fd_sc_hd__clkbuf_1 _5162_ (.A(_2483_),
    .X(_0945_));
 sky130_fd_sc_hd__a22oi_1 _5163_ (.A1(_1549_),
    .A2(\stage_gen[1].mux_gen[13].S.IN1_L5 ),
    .B1(_1550_),
    .B2(\stage_gen[1].mux_gen[13].S.IN1_L3 ),
    .Y(_2484_));
 sky130_fd_sc_hd__o21bai_1 _5164_ (.A1(_2473_),
    .A2(_2484_),
    .B1_N(_0948_),
    .Y(_0947_));
 sky130_fd_sc_hd__a22oi_1 _5165_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[14].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[14].S.IN1_L3 ),
    .Y(_2485_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[7].S.IN1_L1 ),
    .Y(_2486_));
 sky130_fd_sc_hd__o21ai_1 _5167_ (.A1(_2443_),
    .A2(_2485_),
    .B1(_2486_),
    .Y(_0949_));
 sky130_fd_sc_hd__and3_1 _5168_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[7].S.IN1_L2 ),
    .X(_2487_));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(_2487_),
    .X(_0951_));
 sky130_fd_sc_hd__nand2b_1 _5170_ (.A_N(_0951_),
    .B(_2486_),
    .Y(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _5171_ (.A(_2488_),
    .X(_0950_));
 sky130_fd_sc_hd__clkbuf_4 _5172_ (.A(_1369_),
    .X(_2489_));
 sky130_fd_sc_hd__clkbuf_4 _5173_ (.A(_1374_),
    .X(_2490_));
 sky130_fd_sc_hd__a22oi_1 _5174_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[15].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[15].S.IN1_L3 ),
    .Y(_2491_));
 sky130_fd_sc_hd__o21bai_1 _5175_ (.A1(_2473_),
    .A2(_2491_),
    .B1_N(_0953_),
    .Y(_0952_));
 sky130_fd_sc_hd__a22oi_1 _5176_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[16].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[16].S.IN1_L3 ),
    .Y(_2492_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[8].S.IN1_L1 ),
    .Y(_2493_));
 sky130_fd_sc_hd__o21ai_1 _5178_ (.A1(_2443_),
    .A2(_2492_),
    .B1(_2493_),
    .Y(_0954_));
 sky130_fd_sc_hd__and3_1 _5179_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[8].S.IN1_L2 ),
    .X(_2494_));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(_2494_),
    .X(_0956_));
 sky130_fd_sc_hd__nand2b_1 _5181_ (.A_N(_0956_),
    .B(_2493_),
    .Y(_2495_));
 sky130_fd_sc_hd__clkbuf_1 _5182_ (.A(_2495_),
    .X(_0955_));
 sky130_fd_sc_hd__a22oi_1 _5183_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[17].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[17].S.IN1_L3 ),
    .Y(_2496_));
 sky130_fd_sc_hd__o21bai_1 _5184_ (.A1(_2473_),
    .A2(_2496_),
    .B1_N(_0958_),
    .Y(_0957_));
 sky130_fd_sc_hd__a22oi_1 _5185_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[18].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[18].S.IN1_L3 ),
    .Y(_2497_));
 sky130_fd_sc_hd__nand2_1 _5186_ (.A(_2445_),
    .B(\stage_gen[2].mux_gen[9].S.IN1_L1 ),
    .Y(_2498_));
 sky130_fd_sc_hd__o21ai_1 _5187_ (.A1(_2443_),
    .A2(_2497_),
    .B1(_2498_),
    .Y(_0959_));
 sky130_fd_sc_hd__and3_1 _5188_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[9].S.IN1_L2 ),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_1 _5189_ (.A(_2499_),
    .X(_0961_));
 sky130_fd_sc_hd__nand2b_1 _5190_ (.A_N(_0961_),
    .B(_2498_),
    .Y(_2500_));
 sky130_fd_sc_hd__clkbuf_1 _5191_ (.A(_2500_),
    .X(_0960_));
 sky130_fd_sc_hd__a22oi_1 _5192_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[19].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[19].S.IN1_L3 ),
    .Y(_2501_));
 sky130_fd_sc_hd__o21bai_1 _5193_ (.A1(_2473_),
    .A2(_2501_),
    .B1_N(_0963_),
    .Y(_0962_));
 sky130_fd_sc_hd__buf_2 _5194_ (.A(_1421_),
    .X(_2502_));
 sky130_fd_sc_hd__a22oi_1 _5195_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[20].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[20].S.IN1_L3 ),
    .Y(_2503_));
 sky130_fd_sc_hd__buf_2 _5196_ (.A(_1387_),
    .X(_2504_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[10].S.IN1_L1 ),
    .Y(_2505_));
 sky130_fd_sc_hd__o21ai_1 _5198_ (.A1(_2502_),
    .A2(_2503_),
    .B1(_2505_),
    .Y(_0649_));
 sky130_fd_sc_hd__and3_1 _5199_ (.A(_2463_),
    .B(_2452_),
    .C(\stage_gen[2].mux_gen[10].S.IN1_L2 ),
    .X(_2506_));
 sky130_fd_sc_hd__clkbuf_1 _5200_ (.A(_2506_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2b_1 _5201_ (.A_N(_0651_),
    .B(_2505_),
    .Y(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _5202_ (.A(_2507_),
    .X(_0650_));
 sky130_fd_sc_hd__a22oi_1 _5203_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[21].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[21].S.IN1_L3 ),
    .Y(_2508_));
 sky130_fd_sc_hd__o21bai_1 _5204_ (.A1(_2473_),
    .A2(_2508_),
    .B1_N(_0653_),
    .Y(_0652_));
 sky130_fd_sc_hd__a22oi_1 _5205_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[22].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[22].S.IN1_L3 ),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[11].S.IN1_L1 ),
    .Y(_2510_));
 sky130_fd_sc_hd__o21ai_1 _5207_ (.A1(_2502_),
    .A2(_2509_),
    .B1(_2510_),
    .Y(_0654_));
 sky130_fd_sc_hd__buf_2 _5208_ (.A(_1384_),
    .X(_2511_));
 sky130_fd_sc_hd__and3_1 _5209_ (.A(_2463_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[11].S.IN1_L2 ),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _5210_ (.A(_2512_),
    .X(_0656_));
 sky130_fd_sc_hd__nand2b_1 _5211_ (.A_N(_0656_),
    .B(_2510_),
    .Y(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _5212_ (.A(_2513_),
    .X(_0655_));
 sky130_fd_sc_hd__a22oi_1 _5213_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[23].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[23].S.IN1_L3 ),
    .Y(_2514_));
 sky130_fd_sc_hd__o21bai_1 _5214_ (.A1(_2473_),
    .A2(_2514_),
    .B1_N(_0658_),
    .Y(_0657_));
 sky130_fd_sc_hd__a22oi_1 _5215_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[24].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[24].S.IN1_L3 ),
    .Y(_2515_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[12].S.IN1_L1 ),
    .Y(_2516_));
 sky130_fd_sc_hd__o21ai_1 _5217_ (.A1(_2502_),
    .A2(_2515_),
    .B1(_2516_),
    .Y(_0659_));
 sky130_fd_sc_hd__and3_1 _5218_ (.A(_2463_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[12].S.IN1_L2 ),
    .X(_2517_));
 sky130_fd_sc_hd__clkbuf_1 _5219_ (.A(_2517_),
    .X(_0661_));
 sky130_fd_sc_hd__nand2b_1 _5220_ (.A_N(_0661_),
    .B(_2516_),
    .Y(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _5221_ (.A(_2518_),
    .X(_0660_));
 sky130_fd_sc_hd__a22oi_1 _5222_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[25].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[25].S.IN1_L3 ),
    .Y(_2519_));
 sky130_fd_sc_hd__o21bai_1 _5223_ (.A1(_2473_),
    .A2(_2519_),
    .B1_N(_0663_),
    .Y(_0662_));
 sky130_fd_sc_hd__a22oi_1 _5224_ (.A1(_2467_),
    .A2(\stage_gen[1].mux_gen[26].S.IN1_L5 ),
    .B1(_2468_),
    .B2(\stage_gen[1].mux_gen[26].S.IN1_L3 ),
    .Y(_2520_));
 sky130_fd_sc_hd__nand2_1 _5225_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[13].S.IN1_L1 ),
    .Y(_2521_));
 sky130_fd_sc_hd__o21ai_1 _5226_ (.A1(_2502_),
    .A2(_2520_),
    .B1(_2521_),
    .Y(_0664_));
 sky130_fd_sc_hd__buf_2 _5227_ (.A(_1445_),
    .X(_2522_));
 sky130_fd_sc_hd__and3_1 _5228_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[13].S.IN1_L2 ),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_1 _5229_ (.A(_2523_),
    .X(_0666_));
 sky130_fd_sc_hd__nand2b_1 _5230_ (.A_N(_0666_),
    .B(_2521_),
    .Y(_2524_));
 sky130_fd_sc_hd__clkbuf_1 _5231_ (.A(_2524_),
    .X(_0665_));
 sky130_fd_sc_hd__a22oi_1 _5232_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[27].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[27].S.IN1_L3 ),
    .Y(_2525_));
 sky130_fd_sc_hd__o21bai_1 _5233_ (.A1(_2473_),
    .A2(_2525_),
    .B1_N(_0668_),
    .Y(_0667_));
 sky130_fd_sc_hd__clkbuf_4 _5234_ (.A(_1368_),
    .X(_2526_));
 sky130_fd_sc_hd__clkbuf_4 _5235_ (.A(_1373_),
    .X(_2527_));
 sky130_fd_sc_hd__a22oi_1 _5236_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[28].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[28].S.IN1_L3 ),
    .Y(_2528_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[14].S.IN1_L1 ),
    .Y(_2529_));
 sky130_fd_sc_hd__o21ai_1 _5238_ (.A1(_2502_),
    .A2(_2528_),
    .B1(_2529_),
    .Y(_0669_));
 sky130_fd_sc_hd__and3_1 _5239_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[14].S.IN1_L2 ),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_1 _5240_ (.A(_2530_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2b_1 _5241_ (.A_N(_0671_),
    .B(_2529_),
    .Y(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _5242_ (.A(_2531_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_2 _5243_ (.A(_1421_),
    .X(_2532_));
 sky130_fd_sc_hd__a22oi_1 _5244_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[29].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[29].S.IN1_L3 ),
    .Y(_2533_));
 sky130_fd_sc_hd__o21bai_1 _5245_ (.A1(_2532_),
    .A2(_2533_),
    .B1_N(_0673_),
    .Y(_0672_));
 sky130_fd_sc_hd__a22oi_1 _5246_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[30].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[30].S.IN1_L3 ),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[15].S.IN1_L1 ),
    .Y(_2535_));
 sky130_fd_sc_hd__o21ai_1 _5248_ (.A1(_2502_),
    .A2(_2534_),
    .B1(_2535_),
    .Y(_0674_));
 sky130_fd_sc_hd__and3_1 _5249_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[15].S.IN1_L2 ),
    .X(_2536_));
 sky130_fd_sc_hd__clkbuf_1 _5250_ (.A(_2536_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2b_1 _5251_ (.A_N(_0676_),
    .B(_2535_),
    .Y(_2537_));
 sky130_fd_sc_hd__clkbuf_1 _5252_ (.A(_2537_),
    .X(_0675_));
 sky130_fd_sc_hd__a22oi_1 _5253_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[31].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[31].S.IN1_L3 ),
    .Y(_2538_));
 sky130_fd_sc_hd__o21bai_1 _5254_ (.A1(_2532_),
    .A2(_2538_),
    .B1_N(_0678_),
    .Y(_0677_));
 sky130_fd_sc_hd__a22oi_1 _5255_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[32].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[32].S.IN1_L3 ),
    .Y(_2539_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[16].S.IN1_L1 ),
    .Y(_2540_));
 sky130_fd_sc_hd__o21ai_1 _5257_ (.A1(_2502_),
    .A2(_2539_),
    .B1(_2540_),
    .Y(_0679_));
 sky130_fd_sc_hd__and3_1 _5258_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[16].S.IN1_L2 ),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _5259_ (.A(_2541_),
    .X(_0681_));
 sky130_fd_sc_hd__nand2b_1 _5260_ (.A_N(_0681_),
    .B(_2540_),
    .Y(_2542_));
 sky130_fd_sc_hd__clkbuf_1 _5261_ (.A(_2542_),
    .X(_0680_));
 sky130_fd_sc_hd__a22oi_1 _5262_ (.A1(_2489_),
    .A2(\stage_gen[1].mux_gen[33].S.IN1_L5 ),
    .B1(_2490_),
    .B2(\stage_gen[1].mux_gen[33].S.IN1_L3 ),
    .Y(_2543_));
 sky130_fd_sc_hd__o21bai_1 _5263_ (.A1(_2532_),
    .A2(_2543_),
    .B1_N(_0683_),
    .Y(_0682_));
 sky130_fd_sc_hd__a22oi_1 _5264_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[34].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[34].S.IN1_L3 ),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[17].S.IN1_L1 ),
    .Y(_2545_));
 sky130_fd_sc_hd__o21ai_1 _5266_ (.A1(_2502_),
    .A2(_2544_),
    .B1(_2545_),
    .Y(_0684_));
 sky130_fd_sc_hd__and3_1 _5267_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[17].S.IN1_L2 ),
    .X(_2546_));
 sky130_fd_sc_hd__clkbuf_1 _5268_ (.A(_2546_),
    .X(_0686_));
 sky130_fd_sc_hd__nand2b_1 _5269_ (.A_N(_0686_),
    .B(_2545_),
    .Y(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _5270_ (.A(_2547_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_4 _5271_ (.A(_1369_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_4 _5272_ (.A(_1374_),
    .X(_2549_));
 sky130_fd_sc_hd__a22oi_1 _5273_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[35].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[35].S.IN1_L3 ),
    .Y(_2550_));
 sky130_fd_sc_hd__o21bai_1 _5274_ (.A1(_2532_),
    .A2(_2550_),
    .B1_N(_0688_),
    .Y(_0687_));
 sky130_fd_sc_hd__a22oi_1 _5275_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[36].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[36].S.IN1_L3 ),
    .Y(_2551_));
 sky130_fd_sc_hd__nand2_1 _5276_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[18].S.IN1_L1 ),
    .Y(_2552_));
 sky130_fd_sc_hd__o21ai_1 _5277_ (.A1(_2502_),
    .A2(_2551_),
    .B1(_2552_),
    .Y(_0689_));
 sky130_fd_sc_hd__and3_1 _5278_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[18].S.IN1_L2 ),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_1 _5279_ (.A(_2553_),
    .X(_0691_));
 sky130_fd_sc_hd__nand2b_1 _5280_ (.A_N(_0691_),
    .B(_2552_),
    .Y(_2554_));
 sky130_fd_sc_hd__clkbuf_1 _5281_ (.A(_2554_),
    .X(_0690_));
 sky130_fd_sc_hd__a22oi_1 _5282_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[37].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[37].S.IN1_L3 ),
    .Y(_2555_));
 sky130_fd_sc_hd__o21bai_1 _5283_ (.A1(_2532_),
    .A2(_2555_),
    .B1_N(_0693_),
    .Y(_0692_));
 sky130_fd_sc_hd__a22oi_1 _5284_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[38].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[38].S.IN1_L3 ),
    .Y(_2556_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_2504_),
    .B(\stage_gen[2].mux_gen[19].S.IN1_L1 ),
    .Y(_2557_));
 sky130_fd_sc_hd__o21ai_1 _5286_ (.A1(_2502_),
    .A2(_2556_),
    .B1(_2557_),
    .Y(_0694_));
 sky130_fd_sc_hd__and3_1 _5287_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[19].S.IN1_L2 ),
    .X(_2558_));
 sky130_fd_sc_hd__clkbuf_1 _5288_ (.A(_2558_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2b_1 _5289_ (.A_N(_0696_),
    .B(_2557_),
    .Y(_2559_));
 sky130_fd_sc_hd__clkbuf_1 _5290_ (.A(_2559_),
    .X(_0695_));
 sky130_fd_sc_hd__a22oi_1 _5291_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[39].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[39].S.IN1_L3 ),
    .Y(_2560_));
 sky130_fd_sc_hd__o21bai_1 _5292_ (.A1(_2532_),
    .A2(_2560_),
    .B1_N(_0698_),
    .Y(_0697_));
 sky130_fd_sc_hd__clkbuf_4 _5293_ (.A(_1421_),
    .X(_2561_));
 sky130_fd_sc_hd__a22oi_1 _5294_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[40].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[40].S.IN1_L3 ),
    .Y(_2562_));
 sky130_fd_sc_hd__clkbuf_4 _5295_ (.A(_1386_),
    .X(_2563_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[20].S.IN1_L1 ),
    .Y(_2564_));
 sky130_fd_sc_hd__o21ai_1 _5297_ (.A1(_2561_),
    .A2(_2562_),
    .B1(_2564_),
    .Y(_0704_));
 sky130_fd_sc_hd__and3_1 _5298_ (.A(_2522_),
    .B(_2511_),
    .C(\stage_gen[2].mux_gen[20].S.IN1_L2 ),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _5299_ (.A(_2565_),
    .X(_0706_));
 sky130_fd_sc_hd__nand2b_1 _5300_ (.A_N(_0706_),
    .B(_2564_),
    .Y(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _5301_ (.A(_2566_),
    .X(_0705_));
 sky130_fd_sc_hd__a22oi_1 _5302_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[41].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[41].S.IN1_L3 ),
    .Y(_2567_));
 sky130_fd_sc_hd__o21bai_1 _5303_ (.A1(_2532_),
    .A2(_2567_),
    .B1_N(_0708_),
    .Y(_0707_));
 sky130_fd_sc_hd__a22oi_1 _5304_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[42].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[42].S.IN1_L3 ),
    .Y(_2568_));
 sky130_fd_sc_hd__nand2_1 _5305_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[21].S.IN1_L1 ),
    .Y(_2569_));
 sky130_fd_sc_hd__o21ai_1 _5306_ (.A1(_2561_),
    .A2(_2568_),
    .B1(_2569_),
    .Y(_0709_));
 sky130_fd_sc_hd__buf_2 _5307_ (.A(_1384_),
    .X(_2570_));
 sky130_fd_sc_hd__and3_1 _5308_ (.A(_2522_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[21].S.IN1_L2 ),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _5309_ (.A(_2571_),
    .X(_0711_));
 sky130_fd_sc_hd__nand2b_1 _5310_ (.A_N(_0711_),
    .B(_2569_),
    .Y(_2572_));
 sky130_fd_sc_hd__clkbuf_1 _5311_ (.A(_2572_),
    .X(_0710_));
 sky130_fd_sc_hd__a22oi_1 _5312_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[43].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[43].S.IN1_L3 ),
    .Y(_2573_));
 sky130_fd_sc_hd__o21bai_1 _5313_ (.A1(_2532_),
    .A2(_2573_),
    .B1_N(_0713_),
    .Y(_0712_));
 sky130_fd_sc_hd__a22oi_1 _5314_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[44].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[44].S.IN1_L3 ),
    .Y(_2574_));
 sky130_fd_sc_hd__nand2_1 _5315_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[22].S.IN1_L1 ),
    .Y(_2575_));
 sky130_fd_sc_hd__o21ai_1 _5316_ (.A1(_2561_),
    .A2(_2574_),
    .B1(_2575_),
    .Y(_0714_));
 sky130_fd_sc_hd__and3_1 _5317_ (.A(_2522_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[22].S.IN1_L2 ),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _5318_ (.A(_2576_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2b_1 _5319_ (.A_N(_0716_),
    .B(_2575_),
    .Y(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _5320_ (.A(_2577_),
    .X(_0715_));
 sky130_fd_sc_hd__a22oi_1 _5321_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[45].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[45].S.IN1_L3 ),
    .Y(_2578_));
 sky130_fd_sc_hd__o21bai_1 _5322_ (.A1(_2532_),
    .A2(_2578_),
    .B1_N(_0718_),
    .Y(_0717_));
 sky130_fd_sc_hd__a22oi_1 _5323_ (.A1(_2526_),
    .A2(\stage_gen[1].mux_gen[46].S.IN1_L5 ),
    .B1(_2527_),
    .B2(\stage_gen[1].mux_gen[46].S.IN1_L3 ),
    .Y(_2579_));
 sky130_fd_sc_hd__nand2_1 _5324_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[23].S.IN1_L1 ),
    .Y(_2580_));
 sky130_fd_sc_hd__o21ai_1 _5325_ (.A1(_2561_),
    .A2(_2579_),
    .B1(_2580_),
    .Y(_0719_));
 sky130_fd_sc_hd__clkbuf_2 _5326_ (.A(_1445_),
    .X(_2581_));
 sky130_fd_sc_hd__and3_1 _5327_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[23].S.IN1_L2 ),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _5328_ (.A(_2582_),
    .X(_0721_));
 sky130_fd_sc_hd__nand2b_1 _5329_ (.A_N(_0721_),
    .B(_2580_),
    .Y(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _5330_ (.A(_2583_),
    .X(_0720_));
 sky130_fd_sc_hd__a22oi_1 _5331_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[47].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[47].S.IN1_L3 ),
    .Y(_2584_));
 sky130_fd_sc_hd__o21bai_1 _5332_ (.A1(_2532_),
    .A2(_2584_),
    .B1_N(_0723_),
    .Y(_0722_));
 sky130_fd_sc_hd__clkbuf_4 _5333_ (.A(_1368_),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_4 _5334_ (.A(_1373_),
    .X(_2586_));
 sky130_fd_sc_hd__a22oi_1 _5335_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[48].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[48].S.IN1_L3 ),
    .Y(_2587_));
 sky130_fd_sc_hd__nand2_1 _5336_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[24].S.IN1_L1 ),
    .Y(_2588_));
 sky130_fd_sc_hd__o21ai_1 _5337_ (.A1(_2561_),
    .A2(_2587_),
    .B1(_2588_),
    .Y(_0724_));
 sky130_fd_sc_hd__and3_1 _5338_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[24].S.IN1_L2 ),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _5339_ (.A(_2589_),
    .X(_0726_));
 sky130_fd_sc_hd__nand2b_1 _5340_ (.A_N(_0726_),
    .B(_2588_),
    .Y(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _5341_ (.A(_2590_),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _5342_ (.A(_1421_),
    .X(_2591_));
 sky130_fd_sc_hd__a22oi_1 _5343_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[49].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[49].S.IN1_L3 ),
    .Y(_2592_));
 sky130_fd_sc_hd__o21bai_1 _5344_ (.A1(_2591_),
    .A2(_2592_),
    .B1_N(_0728_),
    .Y(_0727_));
 sky130_fd_sc_hd__a22oi_1 _5345_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[50].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[50].S.IN1_L3 ),
    .Y(_2593_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[25].S.IN1_L1 ),
    .Y(_2594_));
 sky130_fd_sc_hd__o21ai_1 _5347_ (.A1(_2561_),
    .A2(_2593_),
    .B1(_2594_),
    .Y(_0729_));
 sky130_fd_sc_hd__and3_1 _5348_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[25].S.IN1_L2 ),
    .X(_2595_));
 sky130_fd_sc_hd__clkbuf_1 _5349_ (.A(_2595_),
    .X(_0731_));
 sky130_fd_sc_hd__nand2b_1 _5350_ (.A_N(_0731_),
    .B(_2594_),
    .Y(_2596_));
 sky130_fd_sc_hd__clkbuf_1 _5351_ (.A(_2596_),
    .X(_0730_));
 sky130_fd_sc_hd__a22oi_1 _5352_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[51].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[51].S.IN1_L3 ),
    .Y(_2597_));
 sky130_fd_sc_hd__o21bai_1 _5353_ (.A1(_2591_),
    .A2(_2597_),
    .B1_N(_0733_),
    .Y(_0732_));
 sky130_fd_sc_hd__a22oi_1 _5354_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[52].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[52].S.IN1_L3 ),
    .Y(_2598_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[26].S.IN1_L1 ),
    .Y(_2599_));
 sky130_fd_sc_hd__o21ai_1 _5356_ (.A1(_2561_),
    .A2(_2598_),
    .B1(_2599_),
    .Y(_0734_));
 sky130_fd_sc_hd__and3_1 _5357_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[26].S.IN1_L2 ),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_1 _5358_ (.A(_2600_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2b_1 _5359_ (.A_N(_0736_),
    .B(_2599_),
    .Y(_2601_));
 sky130_fd_sc_hd__clkbuf_1 _5360_ (.A(_2601_),
    .X(_0735_));
 sky130_fd_sc_hd__a22oi_1 _5361_ (.A1(_2548_),
    .A2(\stage_gen[1].mux_gen[53].S.IN1_L5 ),
    .B1(_2549_),
    .B2(\stage_gen[1].mux_gen[53].S.IN1_L3 ),
    .Y(_2602_));
 sky130_fd_sc_hd__o21bai_1 _5362_ (.A1(_2591_),
    .A2(_2602_),
    .B1_N(_0738_),
    .Y(_0737_));
 sky130_fd_sc_hd__a22oi_1 _5363_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[54].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[54].S.IN1_L3 ),
    .Y(_2603_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[27].S.IN1_L1 ),
    .Y(_2604_));
 sky130_fd_sc_hd__o21ai_1 _5365_ (.A1(_2561_),
    .A2(_2603_),
    .B1(_2604_),
    .Y(_0739_));
 sky130_fd_sc_hd__and3_1 _5366_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[27].S.IN1_L2 ),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _5367_ (.A(_2605_),
    .X(_0741_));
 sky130_fd_sc_hd__nand2b_1 _5368_ (.A_N(_0741_),
    .B(_2604_),
    .Y(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _5369_ (.A(_2606_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_4 _5370_ (.A(_1369_),
    .X(_2607_));
 sky130_fd_sc_hd__buf_4 _5371_ (.A(_1374_),
    .X(_2608_));
 sky130_fd_sc_hd__a22oi_2 _5372_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[55].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[55].S.IN1_L3 ),
    .Y(_2609_));
 sky130_fd_sc_hd__o21bai_1 _5373_ (.A1(_2591_),
    .A2(_2609_),
    .B1_N(_0743_),
    .Y(_0742_));
 sky130_fd_sc_hd__a22oi_1 _5374_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[56].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[56].S.IN1_L3 ),
    .Y(_2610_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[28].S.IN1_L1 ),
    .Y(_2611_));
 sky130_fd_sc_hd__o21ai_1 _5376_ (.A1(_2561_),
    .A2(_2610_),
    .B1(_2611_),
    .Y(_0744_));
 sky130_fd_sc_hd__and3_1 _5377_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[28].S.IN1_L2 ),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _5378_ (.A(_2612_),
    .X(_0746_));
 sky130_fd_sc_hd__nand2b_1 _5379_ (.A_N(_0746_),
    .B(_2611_),
    .Y(_2613_));
 sky130_fd_sc_hd__clkbuf_1 _5380_ (.A(_2613_),
    .X(_0745_));
 sky130_fd_sc_hd__a22oi_1 _5381_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[57].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[57].S.IN1_L3 ),
    .Y(_2614_));
 sky130_fd_sc_hd__o21bai_1 _5382_ (.A1(_2591_),
    .A2(_2614_),
    .B1_N(_0748_),
    .Y(_0747_));
 sky130_fd_sc_hd__a22oi_1 _5383_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[58].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[58].S.IN1_L3 ),
    .Y(_2615_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_2563_),
    .B(\stage_gen[2].mux_gen[29].S.IN1_L1 ),
    .Y(_2616_));
 sky130_fd_sc_hd__o21ai_1 _5385_ (.A1(_2561_),
    .A2(_2615_),
    .B1(_2616_),
    .Y(_0749_));
 sky130_fd_sc_hd__and3_1 _5386_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[29].S.IN1_L2 ),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _5387_ (.A(_2617_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2b_1 _5388_ (.A_N(_0751_),
    .B(_2616_),
    .Y(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _5389_ (.A(_2618_),
    .X(_0750_));
 sky130_fd_sc_hd__a22oi_1 _5390_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[59].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[59].S.IN1_L3 ),
    .Y(_2619_));
 sky130_fd_sc_hd__o21bai_1 _5391_ (.A1(_2591_),
    .A2(_2619_),
    .B1_N(_0753_),
    .Y(_0752_));
 sky130_fd_sc_hd__a22oi_1 _5392_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[60].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[60].S.IN1_L3 ),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[30].S.IN1_L1 ),
    .Y(_2621_));
 sky130_fd_sc_hd__o21ai_1 _5394_ (.A1(_1365_),
    .A2(_2620_),
    .B1(_2621_),
    .Y(_0759_));
 sky130_fd_sc_hd__and3_1 _5395_ (.A(_2581_),
    .B(_2570_),
    .C(\stage_gen[2].mux_gen[30].S.IN1_L2 ),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_1 _5396_ (.A(_2622_),
    .X(_0761_));
 sky130_fd_sc_hd__nand2b_1 _5397_ (.A_N(_0761_),
    .B(_2621_),
    .Y(_2623_));
 sky130_fd_sc_hd__clkbuf_1 _5398_ (.A(_2623_),
    .X(_0760_));
 sky130_fd_sc_hd__a22oi_1 _5399_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[61].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[61].S.IN1_L3 ),
    .Y(_2624_));
 sky130_fd_sc_hd__o21bai_1 _5400_ (.A1(_2591_),
    .A2(_2624_),
    .B1_N(_0763_),
    .Y(_0762_));
 sky130_fd_sc_hd__a22oi_1 _5401_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[62].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[62].S.IN1_L3 ),
    .Y(_2625_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[31].S.IN1_L1 ),
    .Y(_2626_));
 sky130_fd_sc_hd__o21ai_1 _5403_ (.A1(_1365_),
    .A2(_2625_),
    .B1(_2626_),
    .Y(_0764_));
 sky130_fd_sc_hd__and3_1 _5404_ (.A(_2581_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[31].S.IN1_L2 ),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _5405_ (.A(_2627_),
    .X(_0766_));
 sky130_fd_sc_hd__nand2b_1 _5406_ (.A_N(_0766_),
    .B(_2626_),
    .Y(_2628_));
 sky130_fd_sc_hd__clkbuf_1 _5407_ (.A(_2628_),
    .X(_0765_));
 sky130_fd_sc_hd__a22oi_1 _5408_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[63].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[63].S.IN1_L3 ),
    .Y(_2629_));
 sky130_fd_sc_hd__o21bai_1 _5409_ (.A1(_2591_),
    .A2(_2629_),
    .B1_N(_0768_),
    .Y(_0767_));
 sky130_fd_sc_hd__a22oi_1 _5410_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[64].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[64].S.IN1_L3 ),
    .Y(_2630_));
 sky130_fd_sc_hd__nand2_1 _5411_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[32].S.IN1_L1 ),
    .Y(_2631_));
 sky130_fd_sc_hd__o21ai_1 _5412_ (.A1(_1365_),
    .A2(_2630_),
    .B1(_2631_),
    .Y(_0769_));
 sky130_fd_sc_hd__and3_1 _5413_ (.A(_2581_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[32].S.IN1_L2 ),
    .X(_2632_));
 sky130_fd_sc_hd__clkbuf_1 _5414_ (.A(_2632_),
    .X(_0771_));
 sky130_fd_sc_hd__nand2b_1 _5415_ (.A_N(_0771_),
    .B(_2631_),
    .Y(_2633_));
 sky130_fd_sc_hd__clkbuf_1 _5416_ (.A(_2633_),
    .X(_0770_));
 sky130_fd_sc_hd__a22oi_2 _5417_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[65].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[65].S.IN1_L3 ),
    .Y(_2634_));
 sky130_fd_sc_hd__o21bai_1 _5418_ (.A1(_2591_),
    .A2(_2634_),
    .B1_N(_0773_),
    .Y(_0772_));
 sky130_fd_sc_hd__a22oi_1 _5419_ (.A1(_2585_),
    .A2(\stage_gen[1].mux_gen[66].S.IN1_L5 ),
    .B1(_2586_),
    .B2(\stage_gen[1].mux_gen[66].S.IN1_L3 ),
    .Y(_2635_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[33].S.IN1_L1 ),
    .Y(_2636_));
 sky130_fd_sc_hd__o21ai_1 _5421_ (.A1(_1365_),
    .A2(_2635_),
    .B1(_2636_),
    .Y(_0774_));
 sky130_fd_sc_hd__and3_1 _5422_ (.A(_1445_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[33].S.IN1_L2 ),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(_2637_),
    .X(_0776_));
 sky130_fd_sc_hd__or2b_1 _5424_ (.A(_0776_),
    .B_N(_2636_),
    .X(_2638_));
 sky130_fd_sc_hd__clkbuf_1 _5425_ (.A(_2638_),
    .X(_0775_));
 sky130_fd_sc_hd__a22oi_2 _5426_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[67].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[67].S.IN1_L3 ),
    .Y(_2639_));
 sky130_fd_sc_hd__o21bai_1 _5427_ (.A1(_2591_),
    .A2(_2639_),
    .B1_N(_0778_),
    .Y(_0777_));
 sky130_fd_sc_hd__a22oi_1 _5428_ (.A1(_2254_),
    .A2(\stage_gen[1].mux_gen[68].S.IN1_L5 ),
    .B1(_2243_),
    .B2(\stage_gen[1].mux_gen[68].S.IN1_L3 ),
    .Y(_2640_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[34].S.IN1_L1 ),
    .Y(_2641_));
 sky130_fd_sc_hd__o21ai_1 _5430_ (.A1(_1365_),
    .A2(_2640_),
    .B1(_2641_),
    .Y(_0779_));
 sky130_fd_sc_hd__and3_1 _5431_ (.A(_1445_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[34].S.IN1_L2 ),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_1 _5432_ (.A(_2642_),
    .X(_0781_));
 sky130_fd_sc_hd__or2b_1 _5433_ (.A(_0781_),
    .B_N(_2641_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5434_ (.A(_2643_),
    .X(_0780_));
 sky130_fd_sc_hd__a22oi_1 _5435_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[69].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[69].S.IN1_L3 ),
    .Y(_2644_));
 sky130_fd_sc_hd__o21bai_1 _5436_ (.A1(_1380_),
    .A2(_2644_),
    .B1_N(_0783_),
    .Y(_0782_));
 sky130_fd_sc_hd__a22oi_1 _5437_ (.A1(_2254_),
    .A2(\stage_gen[1].mux_gen[70].S.IN1_L5 ),
    .B1(_2243_),
    .B2(\stage_gen[1].mux_gen[70].S.IN1_L3 ),
    .Y(_2645_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[35].S.IN1_L1 ),
    .Y(_2646_));
 sky130_fd_sc_hd__o21ai_1 _5439_ (.A1(_1365_),
    .A2(_2645_),
    .B1(_2646_),
    .Y(_0784_));
 sky130_fd_sc_hd__and3_1 _5440_ (.A(_1445_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[35].S.IN1_L2 ),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2647_),
    .X(_0786_));
 sky130_fd_sc_hd__or2b_1 _5442_ (.A(_0786_),
    .B_N(_2646_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _5443_ (.A(_2648_),
    .X(_0785_));
 sky130_fd_sc_hd__a22oi_1 _5444_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[71].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[71].S.IN1_L3 ),
    .Y(_2649_));
 sky130_fd_sc_hd__o21bai_1 _5445_ (.A1(_1380_),
    .A2(_2649_),
    .B1_N(_0788_),
    .Y(_0787_));
 sky130_fd_sc_hd__a22oi_2 _5446_ (.A1(_2254_),
    .A2(\stage_gen[1].mux_gen[72].S.IN1_L5 ),
    .B1(_2243_),
    .B2(\stage_gen[1].mux_gen[72].S.IN1_L3 ),
    .Y(_2650_));
 sky130_fd_sc_hd__nand2_1 _5447_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[36].S.IN1_L1 ),
    .Y(_2651_));
 sky130_fd_sc_hd__o21ai_1 _5448_ (.A1(_1365_),
    .A2(_2650_),
    .B1(_2651_),
    .Y(_0789_));
 sky130_fd_sc_hd__and3_1 _5449_ (.A(_1445_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[36].S.IN1_L2 ),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5450_ (.A(_2652_),
    .X(_0791_));
 sky130_fd_sc_hd__or2b_1 _5451_ (.A(_0791_),
    .B_N(_2651_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5452_ (.A(_2653_),
    .X(_0790_));
 sky130_fd_sc_hd__a22oi_1 _5453_ (.A1(_2607_),
    .A2(\stage_gen[1].mux_gen[73].S.IN1_L5 ),
    .B1(_2608_),
    .B2(\stage_gen[1].mux_gen[73].S.IN1_L3 ),
    .Y(_2654_));
 sky130_fd_sc_hd__o21bai_1 _5454_ (.A1(_1380_),
    .A2(_2654_),
    .B1_N(_0793_),
    .Y(_0792_));
 sky130_fd_sc_hd__a22oi_1 _5455_ (.A1(_2254_),
    .A2(\stage_gen[1].mux_gen[74].S.IN1_L5 ),
    .B1(_2243_),
    .B2(\stage_gen[1].mux_gen[74].S.IN1_L3 ),
    .Y(_2655_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[37].S.IN1_L1 ),
    .Y(_2656_));
 sky130_fd_sc_hd__o21ai_1 _5457_ (.A1(_1365_),
    .A2(_2655_),
    .B1(_2656_),
    .Y(_0794_));
 sky130_fd_sc_hd__and3_1 _5458_ (.A(_1445_),
    .B(_1361_),
    .C(\stage_gen[2].mux_gen[37].S.IN1_L2 ),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _5459_ (.A(_2657_),
    .X(_0796_));
 sky130_fd_sc_hd__or2b_1 _5460_ (.A(_0796_),
    .B_N(_2656_),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _5461_ (.A(_2658_),
    .X(_0795_));
 sky130_fd_sc_hd__a22oi_1 _5462_ (.A1(_1381_),
    .A2(\stage_gen[1].mux_gen[75].S.IN1_L5 ),
    .B1(_1382_),
    .B2(\stage_gen[1].mux_gen[75].S.IN1_L3 ),
    .Y(_2659_));
 sky130_fd_sc_hd__o21bai_1 _5463_ (.A1(_1380_),
    .A2(_2659_),
    .B1_N(_0798_),
    .Y(_0797_));
 sky130_fd_sc_hd__a22oi_1 _5464_ (.A1(_2254_),
    .A2(\stage_gen[1].mux_gen[76].S.IN1_L5 ),
    .B1(_2243_),
    .B2(\stage_gen[1].mux_gen[76].S.IN1_L3 ),
    .Y(_2660_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_1645_),
    .B(\stage_gen[2].mux_gen[38].S.IN1_L1 ),
    .Y(_2661_));
 sky130_fd_sc_hd__o21ai_1 _5466_ (.A1(_1365_),
    .A2(_2660_),
    .B1(_2661_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2b_1 _5467_ (.A_N(_0801_),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _5468_ (.A(_2662_),
    .X(_0800_));
 sky130_fd_sc_hd__inv_2 _5469_ (.A(\stage_gen[1].genblk1.clks.counter[0] ),
    .Y(_2663_));
 sky130_fd_sc_hd__inv_4 _5470__28 (.A(clknet_1_1__leaf__2236_),
    .Y(net468));
 sky130_fd_sc_hd__inv_4 _5470__29 (.A(clknet_1_1__leaf__2236_),
    .Y(net469));
 sky130_fd_sc_hd__inv_4 _5470__30 (.A(clknet_1_1__leaf__2236_),
    .Y(net470));
 sky130_fd_sc_hd__inv_4 _5470__31 (.A(clknet_1_1__leaf__2236_),
    .Y(net471));
 sky130_fd_sc_hd__inv_4 _5470__32 (.A(clknet_1_0__leaf__2236_),
    .Y(net472));
 sky130_fd_sc_hd__inv_4 _5470__33 (.A(clknet_1_0__leaf__2236_),
    .Y(net473));
 sky130_fd_sc_hd__nand2_2 _5471_ (.A(net461),
    .B(_2663_),
    .Y(_2665_));
 sky130_fd_sc_hd__inv_2 _5472_ (.A(\stage_gen[1].genblk1.clks.counter[9] ),
    .Y(_2666_));
 sky130_fd_sc_hd__inv_2 _5473_ (.A(\stage_gen[1].genblk1.clks.counter[8] ),
    .Y(_2667_));
 sky130_fd_sc_hd__nand2_1 _5474_ (.A(_2666_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__or2_1 _5475_ (.A(\stage_gen[1].genblk1.clks.counter[7] ),
    .B(\stage_gen[1].genblk1.clks.counter[6] ),
    .X(_2669_));
 sky130_fd_sc_hd__nor2_1 _5476_ (.A(_2668_),
    .B(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(\stage_gen[1].genblk1.clks.counter[1] ),
    .B(\stage_gen[1].genblk1.clks.counter[0] ),
    .Y(_2671_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(\stage_gen[1].genblk1.clks.counter[3] ),
    .B(\stage_gen[1].genblk1.clks.counter[2] ),
    .Y(_2672_));
 sky130_fd_sc_hd__nor2_1 _5479_ (.A(_2671_),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_1 _5480_ (.A(\stage_gen[1].genblk1.clks.counter[5] ),
    .B(\stage_gen[1].genblk1.clks.counter[4] ),
    .Y(_2674_));
 sky130_fd_sc_hd__inv_2 _5481_ (.A(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_2673_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_2670_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__o22ai_2 _5484_ (.A1(_2663_),
    .A2(net473),
    .B1(_2665_),
    .B2(_2677_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_2 _5485_ (.A(clknet_1_0__leaf__2017_),
    .B(\stage_gen[1].genblk1.clks.counter[0] ),
    .Y(_2678_));
 sky130_fd_sc_hd__inv_2 _5486__5 (.A(clknet_1_0__leaf__2678_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _5486__6 (.A(clknet_1_1__leaf__2678_),
    .Y(net446));
 sky130_fd_sc_hd__or2_2 _5487_ (.A(\stage_gen[1].genblk1.clks.counter[1] ),
    .B(net446),
    .X(_2680_));
 sky130_fd_sc_hd__nand2_2 _5488_ (.A(net445),
    .B(\stage_gen[1].genblk1.clks.counter[1] ),
    .Y(_2681_));
 sky130_fd_sc_hd__nand2_2 _5489_ (.A(_2680_),
    .B(clknet_1_0__leaf__2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__buf_2 _5490_ (.A(clknet_1_0__leaf__2017_),
    .X(_2683_));
 sky130_fd_sc_hd__nand2_2 _5491_ (.A(_2677_),
    .B(clknet_1_0__leaf__2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand3b_2 _5492_ (.A_N(_2682_),
    .B(clknet_1_0__leaf__2684_),
    .C(_2029_),
    .Y(_2685_));
 sky130_fd_sc_hd__inv_2 _5493__69 (.A(_2685_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _5494_ (.A(\stage_gen[1].genblk1.clks.counter[2] ),
    .Y(_2686_));
 sky130_fd_sc_hd__xor2_2 _5495_ (.A(_2686_),
    .B(clknet_1_1__leaf__2681_),
    .X(_2687_));
 sky130_fd_sc_hd__buf_4 _5496_ (.A(_2019_),
    .X(_2688_));
 sky130_fd_sc_hd__nand3_2 _5497_ (.A(_2687_),
    .B(clknet_1_1__leaf__2684_),
    .C(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__inv_2 _5498__70 (.A(_2689_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _5499_ (.A(\stage_gen[1].genblk1.clks.counter[3] ),
    .Y(_2690_));
 sky130_fd_sc_hd__o21ai_1 _5500_ (.A1(_2686_),
    .A2(_2671_),
    .B1(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__inv_2 _5501_ (.A(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand3b_2 _5502_ (.A_N(_2673_),
    .B(_2670_),
    .C(net460),
    .Y(_2693_));
 sky130_fd_sc_hd__o22ai_2 _5503_ (.A1(_2690_),
    .A2(net472),
    .B1(_2692_),
    .B2(_2693_),
    .Y(_1294_));
 sky130_fd_sc_hd__a21o_2 _5504_ (.A1(_2673_),
    .A2(clknet_1_0__leaf__2017_),
    .B1(\stage_gen[1].genblk1.clks.counter[4] ),
    .X(_2694_));
 sky130_fd_sc_hd__nand3_2 _5505_ (.A(_2673_),
    .B(clknet_1_1__leaf__2683_),
    .C(\stage_gen[1].genblk1.clks.counter[4] ),
    .Y(_2695_));
 sky130_fd_sc_hd__nand2_2 _5506_ (.A(_2694_),
    .B(clknet_1_0__leaf__2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__nand2_2 _5507_ (.A(clknet_1_1__leaf__2684_),
    .B(_2029_),
    .Y(_2697_));
 sky130_fd_sc_hd__nor2_2 _5508_ (.A(_2696_),
    .B(_2697_),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _5509_ (.A(\stage_gen[1].genblk1.clks.counter[5] ),
    .Y(_2698_));
 sky130_fd_sc_hd__nand2_2 _5510_ (.A(clknet_1_1__leaf__2695_),
    .B(_2698_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand3_2 _5511_ (.A(clknet_1_1__leaf__2684_),
    .B(_2688_),
    .C(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__inv_2 _5512__76 (.A(_2700_),
    .Y(net516));
 sky130_fd_sc_hd__nand2_2 _5513_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[1].genblk1.clks.counter[6] ),
    .Y(_2701_));
 sky130_fd_sc_hd__inv_2 _5514__60 (.A(_2701_),
    .Y(net500));
 sky130_fd_sc_hd__nand2_2 _5515_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[1].genblk1.clks.counter[7] ),
    .Y(_2702_));
 sky130_fd_sc_hd__inv_2 _5516__61 (.A(_2702_),
    .Y(net501));
 sky130_fd_sc_hd__buf_1 _5517_ (.A(clknet_1_0__leaf__2017_),
    .X(_2703_));
 sky130_fd_sc_hd__buf_2 _5518_ (.A(_2235_),
    .X(_2704_));
 sky130_fd_sc_hd__or3_4 _5519_ (.A(clknet_1_0__leaf__2703_),
    .B(_2667_),
    .C(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__inv_2 _5520__43 (.A(_2705_),
    .Y(net483));
 sky130_fd_sc_hd__buf_1 _5521_ (.A(clknet_1_0__leaf__2017_),
    .X(_2706_));
 sky130_fd_sc_hd__or3_4 _5522_ (.A(clknet_1_0__leaf__2706_),
    .B(_2666_),
    .C(_2704_),
    .X(_2707_));
 sky130_fd_sc_hd__inv_2 _5523__48 (.A(_2707_),
    .Y(net488));
 sky130_fd_sc_hd__nand2_2 _5524_ (.A(clknet_1_0__leaf__2684_),
    .B(_2034_),
    .Y(_2708_));
 sky130_fd_sc_hd__nand3_2 _5525_ (.A(_2677_),
    .B(clknet_1_0__leaf__2018_),
    .C(_2240_),
    .Y(_2709_));
 sky130_fd_sc_hd__nand3_2 _5526_ (.A(_2708_),
    .B(_2688_),
    .C(_2709_),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _5527_ (.A(\stage_gen[2].genblk1.clks.counter[9] ),
    .Y(_2710_));
 sky130_fd_sc_hd__inv_2 _5528_ (.A(\stage_gen[2].genblk1.clks.counter[8] ),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_1 _5529_ (.A(_2710_),
    .B(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__nor2_1 _5530_ (.A(\stage_gen[2].genblk1.clks.counter[7] ),
    .B(\stage_gen[2].genblk1.clks.counter[5] ),
    .Y(_2713_));
 sky130_fd_sc_hd__inv_2 _5531_ (.A(\stage_gen[2].genblk1.clks.counter[6] ),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_2713_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__nor2_1 _5533_ (.A(_2712_),
    .B(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(\stage_gen[2].genblk1.clks.counter[1] ),
    .B(\stage_gen[2].genblk1.clks.counter[0] ),
    .Y(_2717_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(\stage_gen[2].genblk1.clks.counter[3] ),
    .B(\stage_gen[2].genblk1.clks.counter[2] ),
    .Y(_2718_));
 sky130_fd_sc_hd__nor2_1 _5536_ (.A(_2717_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_1 _5537_ (.A(_2719_),
    .B(\stage_gen[2].genblk1.clks.counter[4] ),
    .Y(_2720_));
 sky130_fd_sc_hd__nand3_2 _5538_ (.A(_2716_),
    .B(_2720_),
    .C(net459),
    .Y(_2721_));
 sky130_fd_sc_hd__inv_2 _5539_ (.A(\stage_gen[2].genblk1.clks.counter[0] ),
    .Y(_2722_));
 sky130_fd_sc_hd__nor2_2 _5540_ (.A(_2722_),
    .B(clknet_1_0__leaf__2236_),
    .Y(_2723_));
 sky130_fd_sc_hd__a21oi_2 _5541_ (.A1(clknet_1_1__leaf__2721_),
    .A2(_2722_),
    .B1(_2723_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_2 _5542_ (.A(clknet_3_4__leaf_CLK),
    .B(\stage_gen[2].genblk1.clks.counter[0] ),
    .Y(_2724_));
 sky130_fd_sc_hd__inv_2 _5543__7 (.A(clknet_1_0__leaf__2724_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _5543__8 (.A(clknet_1_1__leaf__2724_),
    .Y(net448));
 sky130_fd_sc_hd__or2_2 _5544_ (.A(\stage_gen[2].genblk1.clks.counter[1] ),
    .B(net448),
    .X(_2726_));
 sky130_fd_sc_hd__nand2_2 _5545_ (.A(net447),
    .B(\stage_gen[2].genblk1.clks.counter[1] ),
    .Y(_2727_));
 sky130_fd_sc_hd__nand2_2 _5546_ (.A(_2726_),
    .B(clknet_1_1__leaf__2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(_2716_),
    .B(_2720_),
    .Y(_2729_));
 sky130_fd_sc_hd__nand2_2 _5548_ (.A(_2729_),
    .B(clknet_1_0__leaf__2683_),
    .Y(_2730_));
 sky130_fd_sc_hd__nand3b_2 _5549_ (.A_N(_2728_),
    .B(clknet_1_1__leaf__2730_),
    .C(_2029_),
    .Y(_2731_));
 sky130_fd_sc_hd__inv_2 _5550__71 (.A(_2731_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _5551_ (.A(\stage_gen[2].genblk1.clks.counter[2] ),
    .Y(_2732_));
 sky130_fd_sc_hd__xor2_2 _5552_ (.A(_2732_),
    .B(clknet_1_0__leaf__2727_),
    .X(_2733_));
 sky130_fd_sc_hd__nand3_2 _5553_ (.A(_2733_),
    .B(clknet_1_1__leaf__2730_),
    .C(_2688_),
    .Y(_2734_));
 sky130_fd_sc_hd__inv_2 _5554__72 (.A(_2734_),
    .Y(net512));
 sky130_fd_sc_hd__nor2_1 _5555_ (.A(_2732_),
    .B(_2717_),
    .Y(_2735_));
 sky130_fd_sc_hd__xnor2_1 _5556_ (.A(\stage_gen[2].genblk1.clks.counter[3] ),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__nand2_2 _5557_ (.A(clknet_1_0__leaf__2236_),
    .B(\stage_gen[2].genblk1.clks.counter[3] ),
    .Y(_2737_));
 sky130_fd_sc_hd__o21ai_2 _5558_ (.A1(_2736_),
    .A2(clknet_1_0__leaf__2721_),
    .B1(_2737_),
    .Y(_1305_));
 sky130_fd_sc_hd__a21o_2 _5559_ (.A1(_2719_),
    .A2(clknet_1_0__leaf__2683_),
    .B1(\stage_gen[2].genblk1.clks.counter[4] ),
    .X(_2738_));
 sky130_fd_sc_hd__nand3_2 _5560_ (.A(clknet_1_0__leaf__2730_),
    .B(_2738_),
    .C(_2688_),
    .Y(_2739_));
 sky130_fd_sc_hd__inv_2 _5561__77 (.A(_2739_),
    .Y(net517));
 sky130_fd_sc_hd__nand2_2 _5562_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[2].genblk1.clks.counter[5] ),
    .Y(_2740_));
 sky130_fd_sc_hd__inv_2 _5563__62 (.A(_2740_),
    .Y(net502));
 sky130_fd_sc_hd__or3_4 _5564_ (.A(clknet_1_0__leaf__2706_),
    .B(_2714_),
    .C(_2704_),
    .X(_2741_));
 sky130_fd_sc_hd__inv_2 _5565__49 (.A(_2741_),
    .Y(net489));
 sky130_fd_sc_hd__nand2_2 _5566_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[2].genblk1.clks.counter[7] ),
    .Y(_2742_));
 sky130_fd_sc_hd__inv_2 _5567__63 (.A(_2742_),
    .Y(net503));
 sky130_fd_sc_hd__or3_4 _5568_ (.A(clknet_1_0__leaf__2706_),
    .B(_2711_),
    .C(_2704_),
    .X(_2743_));
 sky130_fd_sc_hd__inv_2 _5569__50 (.A(_2743_),
    .Y(net490));
 sky130_fd_sc_hd__or3_4 _5570_ (.A(clknet_1_0__leaf__2706_),
    .B(_2710_),
    .C(_2704_),
    .X(_2744_));
 sky130_fd_sc_hd__inv_2 _5571__51 (.A(_2744_),
    .Y(net491));
 sky130_fd_sc_hd__nand2_2 _5572_ (.A(clknet_1_0__leaf__2730_),
    .B(_1380_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand3_2 _5573_ (.A(_2729_),
    .B(clknet_1_0__leaf__2018_),
    .C(_1359_),
    .Y(_2746_));
 sky130_fd_sc_hd__nand3_2 _5574_ (.A(_2745_),
    .B(_2688_),
    .C(_2746_),
    .Y(_1312_));
 sky130_fd_sc_hd__inv_2 _5575_ (.A(\stage_gen[3].genblk1.clks.counter[0] ),
    .Y(_2747_));
 sky130_fd_sc_hd__nand2_2 _5576_ (.A(net458),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__inv_2 _5577_ (.A(\stage_gen[3].genblk1.clks.counter[7] ),
    .Y(_2749_));
 sky130_fd_sc_hd__inv_2 _5578_ (.A(\stage_gen[3].genblk1.clks.counter[6] ),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_2749_),
    .B(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(\stage_gen[3].genblk1.clks.counter[5] ),
    .Y(_2752_));
 sky130_fd_sc_hd__inv_2 _5581_ (.A(\stage_gen[3].genblk1.clks.counter[4] ),
    .Y(_2753_));
 sky130_fd_sc_hd__nand2_1 _5582_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nor2_1 _5583_ (.A(_2751_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(\stage_gen[3].genblk1.clks.counter[9] ),
    .B(\stage_gen[3].genblk1.clks.counter[8] ),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(\stage_gen[3].genblk1.clks.counter[1] ),
    .B(\stage_gen[3].genblk1.clks.counter[0] ),
    .Y(_2757_));
 sky130_fd_sc_hd__inv_2 _5586_ (.A(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(\stage_gen[3].genblk1.clks.counter[3] ),
    .B(\stage_gen[3].genblk1.clks.counter[2] ),
    .Y(_2759_));
 sky130_fd_sc_hd__inv_2 _5588_ (.A(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__nand2_1 _5589_ (.A(_2758_),
    .B(_2760_),
    .Y(_2761_));
 sky130_fd_sc_hd__nand3_2 _5590_ (.A(_2755_),
    .B(_2756_),
    .C(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__o22ai_2 _5591_ (.A1(_2747_),
    .A2(net471),
    .B1(_2748_),
    .B2(_2762_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_2 _5592_ (.A(clknet_3_4__leaf_CLK),
    .B(\stage_gen[3].genblk1.clks.counter[0] ),
    .Y(_2763_));
 sky130_fd_sc_hd__inv_2 _5593__10 (.A(clknet_1_1__leaf__2763_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _5593__9 (.A(clknet_1_0__leaf__2763_),
    .Y(net449));
 sky130_fd_sc_hd__or2_2 _5594_ (.A(\stage_gen[3].genblk1.clks.counter[1] ),
    .B(net450),
    .X(_2765_));
 sky130_fd_sc_hd__nand2_2 _5595_ (.A(net449),
    .B(\stage_gen[3].genblk1.clks.counter[1] ),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_2 _5596_ (.A(_2765_),
    .B(clknet_1_0__leaf__2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__nand2_2 _5597_ (.A(_2762_),
    .B(clknet_1_0__leaf__2683_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand3b_2 _5598_ (.A_N(_2767_),
    .B(clknet_1_0__leaf__2768_),
    .C(_2029_),
    .Y(_2769_));
 sky130_fd_sc_hd__inv_2 _5599__73 (.A(_2769_),
    .Y(net513));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(_2758_),
    .B(\stage_gen[3].genblk1.clks.counter[2] ),
    .Y(_2770_));
 sky130_fd_sc_hd__inv_2 _5601_ (.A(\stage_gen[3].genblk1.clks.counter[2] ),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_2 _5602_ (.A(clknet_1_1__leaf__2766_),
    .B(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__o21ai_2 _5603_ (.A1(net442),
    .A2(_2770_),
    .B1(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__inv_2 _5604__59 (.A(_2773_),
    .Y(net499));
 sky130_fd_sc_hd__nand3_2 _5605_ (.A(net499),
    .B(clknet_1_1__leaf__2768_),
    .C(_2029_),
    .Y(_2775_));
 sky130_fd_sc_hd__inv_2 _5606__78 (.A(_2775_),
    .Y(net518));
 sky130_fd_sc_hd__o21ba_2 _5607_ (.A1(net441),
    .A2(_2770_),
    .B1_N(\stage_gen[3].genblk1.clks.counter[3] ),
    .X(_2776_));
 sky130_fd_sc_hd__nand2_2 _5608_ (.A(clknet_1_1__leaf__2768_),
    .B(_2029_),
    .Y(_2777_));
 sky130_fd_sc_hd__nor2_2 _5609_ (.A(_2776_),
    .B(_2777_),
    .Y(_1316_));
 sky130_fd_sc_hd__or3_4 _5610_ (.A(clknet_1_0__leaf__2706_),
    .B(_2753_),
    .C(_2704_),
    .X(_2778_));
 sky130_fd_sc_hd__inv_2 _5611__52 (.A(_2778_),
    .Y(net492));
 sky130_fd_sc_hd__nand2_2 _5612_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[3].genblk1.clks.counter[5] ),
    .Y(_2779_));
 sky130_fd_sc_hd__inv_2 _5613__64 (.A(_2779_),
    .Y(net504));
 sky130_fd_sc_hd__or3_4 _5614_ (.A(clknet_1_0__leaf__2706_),
    .B(_2750_),
    .C(_2704_),
    .X(_2780_));
 sky130_fd_sc_hd__inv_2 _5615__53 (.A(_2780_),
    .Y(net493));
 sky130_fd_sc_hd__nand2_2 _5616_ (.A(clknet_1_0__leaf__1290_),
    .B(\stage_gen[3].genblk1.clks.counter[7] ),
    .Y(_2781_));
 sky130_fd_sc_hd__inv_2 _5617__65 (.A(_2781_),
    .Y(net505));
 sky130_fd_sc_hd__buf_6 _5618_ (.A(_2235_),
    .X(_2782_));
 sky130_fd_sc_hd__or3b_4 _5619_ (.A(clknet_1_1__leaf__2683_),
    .B(_2782_),
    .C_N(\stage_gen[3].genblk1.clks.counter[8] ),
    .X(_2783_));
 sky130_fd_sc_hd__inv_2 _5620__39 (.A(_2783_),
    .Y(net479));
 sky130_fd_sc_hd__or3b_4 _5621_ (.A(clknet_1_1__leaf__2683_),
    .B(_2782_),
    .C_N(\stage_gen[3].genblk1.clks.counter[9] ),
    .X(_2784_));
 sky130_fd_sc_hd__inv_2 _5622__40 (.A(_2784_),
    .Y(net480));
 sky130_fd_sc_hd__nand2_2 _5623_ (.A(clknet_1_0__leaf__2768_),
    .B(_1566_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand3_2 _5624_ (.A(_2762_),
    .B(clknet_1_0__leaf__2018_),
    .C(_1579_),
    .Y(_2786_));
 sky130_fd_sc_hd__nand3_2 _5625_ (.A(_2785_),
    .B(_2688_),
    .C(_2786_),
    .Y(_1323_));
 sky130_fd_sc_hd__inv_2 _5626_ (.A(\stage_gen[4].genblk1.clks.counter[0] ),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2_2 _5627_ (.A(net457),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__inv_2 _5628_ (.A(\stage_gen[4].genblk1.clks.counter[2] ),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(\stage_gen[4].genblk1.clks.counter[1] ),
    .B(\stage_gen[4].genblk1.clks.counter[0] ),
    .Y(_2790_));
 sky130_fd_sc_hd__nor2_1 _5630_ (.A(_2789_),
    .B(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__nor2_1 _5631_ (.A(\stage_gen[4].genblk1.clks.counter[8] ),
    .B(\stage_gen[4].genblk1.clks.counter[7] ),
    .Y(_2792_));
 sky130_fd_sc_hd__inv_2 _5632_ (.A(\stage_gen[4].genblk1.clks.counter[4] ),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_2792_),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__nor2_1 _5634_ (.A(_2791_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__nor2_1 _5635_ (.A(\stage_gen[4].genblk1.clks.counter[5] ),
    .B(\stage_gen[4].genblk1.clks.counter[3] ),
    .Y(_2796_));
 sky130_fd_sc_hd__nor2_1 _5636_ (.A(\stage_gen[4].genblk1.clks.counter[9] ),
    .B(\stage_gen[4].genblk1.clks.counter[6] ),
    .Y(_2797_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(_2796_),
    .B(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2_1 _5638_ (.A(_2795_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__o22ai_2 _5639_ (.A1(_2787_),
    .A2(net470),
    .B1(_2788_),
    .B2(_2799_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_2 _5640_ (.A(clknet_3_5__leaf_CLK),
    .B(\stage_gen[4].genblk1.clks.counter[0] ),
    .Y(_2800_));
 sky130_fd_sc_hd__inv_2 _5641__11 (.A(clknet_1_1__leaf__2800_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _5641__12 (.A(clknet_1_0__leaf__2800_),
    .Y(net452));
 sky130_fd_sc_hd__or2_2 _5642_ (.A(\stage_gen[4].genblk1.clks.counter[1] ),
    .B(net452),
    .X(_2802_));
 sky130_fd_sc_hd__nand2_2 _5643_ (.A(net451),
    .B(\stage_gen[4].genblk1.clks.counter[1] ),
    .Y(_2803_));
 sky130_fd_sc_hd__nand2_2 _5644_ (.A(_2802_),
    .B(clknet_1_1__leaf__2803_),
    .Y(_2804_));
 sky130_fd_sc_hd__nand2_2 _5645_ (.A(_2799_),
    .B(clknet_1_1__leaf__2018_),
    .Y(_2805_));
 sky130_fd_sc_hd__nand3b_2 _5646_ (.A_N(_2804_),
    .B(clknet_1_0__leaf__2805_),
    .C(_2029_),
    .Y(_2806_));
 sky130_fd_sc_hd__inv_2 _5647__74 (.A(_2806_),
    .Y(net514));
 sky130_fd_sc_hd__xor2_2 _5648_ (.A(_2789_),
    .B(clknet_1_0__leaf__2803_),
    .X(_2807_));
 sky130_fd_sc_hd__nand3_2 _5649_ (.A(clknet_1_1__leaf__2805_),
    .B(_2807_),
    .C(_2029_),
    .Y(_2808_));
 sky130_fd_sc_hd__inv_2 _5650__75 (.A(_2808_),
    .Y(net515));
 sky130_fd_sc_hd__nand2_2 _5651_ (.A(clknet_1_1__leaf__1290_),
    .B(\stage_gen[4].genblk1.clks.counter[3] ),
    .Y(_2809_));
 sky130_fd_sc_hd__inv_2 _5652__66 (.A(_2809_),
    .Y(net506));
 sky130_fd_sc_hd__or3_4 _5653_ (.A(clknet_1_1__leaf__2706_),
    .B(_2793_),
    .C(_2704_),
    .X(_2810_));
 sky130_fd_sc_hd__inv_2 _5654__54 (.A(_2810_),
    .Y(net494));
 sky130_fd_sc_hd__nand2_2 _5655_ (.A(clknet_1_1__leaf__1290_),
    .B(\stage_gen[4].genblk1.clks.counter[5] ),
    .Y(_2811_));
 sky130_fd_sc_hd__inv_2 _5656__67 (.A(_2811_),
    .Y(net507));
 sky130_fd_sc_hd__or3b_4 _5657_ (.A(clknet_1_1__leaf__2683_),
    .B(_2782_),
    .C_N(\stage_gen[4].genblk1.clks.counter[6] ),
    .X(_2812_));
 sky130_fd_sc_hd__inv_2 _5658__41 (.A(_2812_),
    .Y(net481));
 sky130_fd_sc_hd__nand2_2 _5659_ (.A(clknet_1_1__leaf__1290_),
    .B(\stage_gen[4].genblk1.clks.counter[7] ),
    .Y(_2813_));
 sky130_fd_sc_hd__inv_2 _5660__68 (.A(_2813_),
    .Y(net508));
 sky130_fd_sc_hd__or3b_4 _5661_ (.A(clknet_1_1__leaf__2683_),
    .B(_2782_),
    .C_N(\stage_gen[4].genblk1.clks.counter[8] ),
    .X(_2814_));
 sky130_fd_sc_hd__inv_2 _5662__42 (.A(_2814_),
    .Y(net482));
 sky130_fd_sc_hd__or3b_4 _5663_ (.A(clknet_1_1__leaf__2703_),
    .B(_2782_),
    .C_N(\stage_gen[4].genblk1.clks.counter[9] ),
    .X(_2815_));
 sky130_fd_sc_hd__inv_2 _5664__44 (.A(_2815_),
    .Y(net484));
 sky130_fd_sc_hd__nand2_2 _5665_ (.A(clknet_1_0__leaf__2805_),
    .B(_1799_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand3_2 _5666_ (.A(_2799_),
    .B(clknet_1_1__leaf__2018_),
    .C(_1811_),
    .Y(_2817_));
 sky130_fd_sc_hd__nand3_2 _5667_ (.A(_2816_),
    .B(_2688_),
    .C(_2817_),
    .Y(_1334_));
 sky130_fd_sc_hd__inv_2 _5668_ (.A(\stage_gen[5].genblk1.clks.counter[0] ),
    .Y(_2818_));
 sky130_fd_sc_hd__nand2_2 _5669_ (.A(net456),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(\stage_gen[5].genblk1.clks.counter[1] ),
    .B(\stage_gen[5].genblk1.clks.counter[0] ),
    .Y(_2820_));
 sky130_fd_sc_hd__inv_2 _5671_ (.A(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__nor2_1 _5672_ (.A(\stage_gen[5].genblk1.clks.counter[9] ),
    .B(\stage_gen[5].genblk1.clks.counter[8] ),
    .Y(_2822_));
 sky130_fd_sc_hd__nor2_1 _5673_ (.A(\stage_gen[5].genblk1.clks.counter[7] ),
    .B(\stage_gen[5].genblk1.clks.counter[6] ),
    .Y(_2823_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_2822_),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__nor2_1 _5675_ (.A(_2821_),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__nor2_1 _5676_ (.A(\stage_gen[5].genblk1.clks.counter[5] ),
    .B(\stage_gen[5].genblk1.clks.counter[4] ),
    .Y(_2826_));
 sky130_fd_sc_hd__nor2_1 _5677_ (.A(\stage_gen[5].genblk1.clks.counter[3] ),
    .B(\stage_gen[5].genblk1.clks.counter[2] ),
    .Y(_2827_));
 sky130_fd_sc_hd__and2_1 _5678_ (.A(_2826_),
    .B(_2827_),
    .X(_2828_));
 sky130_fd_sc_hd__nand2_2 _5679_ (.A(_2825_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__o22ai_2 _5680_ (.A1(_2818_),
    .A2(net469),
    .B1(_2819_),
    .B2(_2829_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_2 _5681_ (.A(_2829_),
    .B(clknet_1_1__leaf__2018_),
    .Y(_2830_));
 sky130_fd_sc_hd__nand3_2 _5682_ (.A(clknet_1_1__leaf__2830_),
    .B(\stage_gen[5].genblk1.clks.counter[1] ),
    .C(_2029_),
    .Y(_2831_));
 sky130_fd_sc_hd__nor2_2 _5683_ (.A(clknet_1_1__leaf__2022_),
    .B(_2829_),
    .Y(_2832_));
 sky130_fd_sc_hd__nand2_2 _5684_ (.A(_2832_),
    .B(\stage_gen[5].genblk1.clks.counter[0] ),
    .Y(_2833_));
 sky130_fd_sc_hd__nand2_2 _5685_ (.A(_2831_),
    .B(_2833_),
    .Y(_1336_));
 sky130_fd_sc_hd__or3b_4 _5686_ (.A(clknet_1_1__leaf__2703_),
    .B(_2782_),
    .C_N(\stage_gen[5].genblk1.clks.counter[2] ),
    .X(_2834_));
 sky130_fd_sc_hd__inv_2 _5687__45 (.A(_2834_),
    .Y(net485));
 sky130_fd_sc_hd__or3b_4 _5688_ (.A(clknet_1_1__leaf__2703_),
    .B(_2782_),
    .C_N(\stage_gen[5].genblk1.clks.counter[3] ),
    .X(_2835_));
 sky130_fd_sc_hd__inv_2 _5689__46 (.A(_2835_),
    .Y(net486));
 sky130_fd_sc_hd__or3b_4 _5690_ (.A(clknet_1_1__leaf__2703_),
    .B(_2782_),
    .C_N(\stage_gen[5].genblk1.clks.counter[4] ),
    .X(_2836_));
 sky130_fd_sc_hd__inv_2 _5691__47 (.A(_2836_),
    .Y(net487));
 sky130_fd_sc_hd__nand2_2 _5692_ (.A(clknet_1_1__leaf__2236_),
    .B(\stage_gen[5].genblk1.clks.counter[5] ),
    .Y(_2837_));
 sky130_fd_sc_hd__inv_2 _5693__34 (.A(_2837_),
    .Y(net474));
 sky130_fd_sc_hd__or3b_2 _5694_ (.A(clknet_1_0__leaf__2703_),
    .B(_2235_),
    .C_N(\stage_gen[5].genblk1.clks.counter[6] ),
    .X(_2838_));
 sky130_fd_sc_hd__inv_2 _5695__23 (.A(_2838_),
    .Y(net463));
 sky130_fd_sc_hd__nand2_2 _5696_ (.A(clknet_1_1__leaf__2236_),
    .B(\stage_gen[5].genblk1.clks.counter[7] ),
    .Y(_2839_));
 sky130_fd_sc_hd__inv_2 _5697__35 (.A(_2839_),
    .Y(net475));
 sky130_fd_sc_hd__or3b_2 _5698_ (.A(clknet_1_1__leaf__2703_),
    .B(_2235_),
    .C_N(\stage_gen[5].genblk1.clks.counter[8] ),
    .X(_2840_));
 sky130_fd_sc_hd__inv_2 _5699__24 (.A(_2840_),
    .Y(net464));
 sky130_fd_sc_hd__or3b_2 _5700_ (.A(clknet_1_1__leaf__2703_),
    .B(_2235_),
    .C_N(\stage_gen[5].genblk1.clks.counter[9] ),
    .X(_2841_));
 sky130_fd_sc_hd__inv_2 _5701__25 (.A(_2841_),
    .Y(net465));
 sky130_fd_sc_hd__nand2_2 _5702_ (.A(clknet_1_0__leaf__2830_),
    .B(_1917_),
    .Y(_2842_));
 sky130_fd_sc_hd__nand3_2 _5703_ (.A(_2829_),
    .B(clknet_1_1__leaf__2018_),
    .C(_1924_),
    .Y(_2843_));
 sky130_fd_sc_hd__nand3_2 _5704_ (.A(_2842_),
    .B(_2688_),
    .C(_2843_),
    .Y(_1345_));
 sky130_fd_sc_hd__nor2_2 _5705_ (.A(clknet_1_0__leaf__2018_),
    .B(\stage_gen[6].genblk1.clks.counter[0] ),
    .Y(_2844_));
 sky130_fd_sc_hd__inv_2 _5706_ (.A(\stage_gen[6].genblk1.clks.counter[9] ),
    .Y(_2845_));
 sky130_fd_sc_hd__inv_2 _5707_ (.A(\stage_gen[6].genblk1.clks.counter[8] ),
    .Y(_2846_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_2845_),
    .B(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _5709_ (.A(\stage_gen[6].genblk1.clks.counter[7] ),
    .B(\stage_gen[6].genblk1.clks.counter[6] ),
    .Y(_2848_));
 sky130_fd_sc_hd__nor2_1 _5710_ (.A(\stage_gen[6].genblk1.clks.counter[5] ),
    .B(\stage_gen[6].genblk1.clks.counter[4] ),
    .Y(_2849_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_2848_),
    .B(_2849_),
    .Y(_2850_));
 sky130_fd_sc_hd__nor2_1 _5712_ (.A(_2847_),
    .B(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__inv_2 _5713_ (.A(\stage_gen[6].genblk1.clks.counter[2] ),
    .Y(_2852_));
 sky130_fd_sc_hd__inv_2 _5714_ (.A(\stage_gen[6].genblk1.clks.counter[1] ),
    .Y(_2853_));
 sky130_fd_sc_hd__nand2_1 _5715_ (.A(_2852_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__or2_1 _5716_ (.A(\stage_gen[6].genblk1.clks.counter[3] ),
    .B(\stage_gen[6].genblk1.clks.counter[0] ),
    .X(_2855_));
 sky130_fd_sc_hd__nor2_1 _5717_ (.A(_2854_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(_2851_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__nand2_2 _5719_ (.A(_2857_),
    .B(clknet_1_1__leaf__2683_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand2_2 _5720_ (.A(clknet_1_0__leaf__2858_),
    .B(_2019_),
    .Y(_2859_));
 sky130_fd_sc_hd__nor2_2 _5721_ (.A(_2844_),
    .B(_2859_),
    .Y(_1346_));
 sky130_fd_sc_hd__or3_4 _5722_ (.A(clknet_1_1__leaf__2706_),
    .B(_2853_),
    .C(_2704_),
    .X(_2860_));
 sky130_fd_sc_hd__inv_2 _5723__55 (.A(_2860_),
    .Y(net495));
 sky130_fd_sc_hd__or3_4 _5724_ (.A(clknet_1_1__leaf__2706_),
    .B(_2852_),
    .C(_2704_),
    .X(_2861_));
 sky130_fd_sc_hd__inv_2 _5725__56 (.A(_2861_),
    .Y(net496));
 sky130_fd_sc_hd__nand2_2 _5726_ (.A(clknet_1_0__leaf__2236_),
    .B(\stage_gen[6].genblk1.clks.counter[3] ),
    .Y(_2862_));
 sky130_fd_sc_hd__inv_2 _5727__36 (.A(_2862_),
    .Y(net476));
 sky130_fd_sc_hd__or3b_2 _5728_ (.A(clknet_1_0__leaf__2703_),
    .B(_2235_),
    .C_N(\stage_gen[6].genblk1.clks.counter[4] ),
    .X(_2863_));
 sky130_fd_sc_hd__inv_2 _5729__26 (.A(_2863_),
    .Y(net466));
 sky130_fd_sc_hd__nand2_2 _5730_ (.A(clknet_1_0__leaf__2236_),
    .B(\stage_gen[6].genblk1.clks.counter[5] ),
    .Y(_2864_));
 sky130_fd_sc_hd__inv_2 _5731__37 (.A(_2864_),
    .Y(net477));
 sky130_fd_sc_hd__or3b_2 _5732_ (.A(clknet_1_0__leaf__2703_),
    .B(_2235_),
    .C_N(\stage_gen[6].genblk1.clks.counter[6] ),
    .X(_2865_));
 sky130_fd_sc_hd__inv_2 _5733__27 (.A(_2865_),
    .Y(net467));
 sky130_fd_sc_hd__nand2_2 _5734_ (.A(clknet_1_0__leaf__2236_),
    .B(\stage_gen[6].genblk1.clks.counter[7] ),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _5735__38 (.A(_2866_),
    .Y(net478));
 sky130_fd_sc_hd__or3_4 _5736_ (.A(clknet_1_1__leaf__2706_),
    .B(_2846_),
    .C(_2782_),
    .X(_2867_));
 sky130_fd_sc_hd__inv_2 _5737__57 (.A(_2867_),
    .Y(net497));
 sky130_fd_sc_hd__or3_4 _5738_ (.A(clknet_1_1__leaf__2017_),
    .B(_2845_),
    .C(_2782_),
    .X(_2868_));
 sky130_fd_sc_hd__inv_2 _5739__58 (.A(_2868_),
    .Y(net498));
 sky130_fd_sc_hd__nand2_2 _5740_ (.A(clknet_1_1__leaf__2858_),
    .B(_1973_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand3_2 _5741_ (.A(_2857_),
    .B(clknet_1_1__leaf__2018_),
    .C(_1978_),
    .Y(_2870_));
 sky130_fd_sc_hd__nand3_2 _5742_ (.A(_2869_),
    .B(_2688_),
    .C(_2870_),
    .Y(_1356_));
 sky130_fd_sc_hd__mux2_2 _5743_ (.A0(net468),
    .A1(clknet_1_1__leaf__2022_),
    .S(_2001_),
    .X(_2871_));
 sky130_fd_sc_hd__buf_6 _5744_ (.A(_2871_),
    .X(_1357_));
 sky130_fd_sc_hd__dfxtp_1 _5745_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_1291_),
    .Q(\stage_gen[1].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5746_ (.CLK(clknet_3_0__leaf_CLK),
    .D(net509),
    .Q(\stage_gen[1].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5747_ (.CLK(clknet_3_0__leaf_CLK),
    .D(net510),
    .Q(\stage_gen[1].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5748_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_1294_),
    .Q(\stage_gen[1].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5749_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_1295_),
    .Q(\stage_gen[1].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5750_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net516),
    .Q(\stage_gen[1].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5751_ (.CLK(clknet_3_0__leaf_CLK),
    .D(net500),
    .Q(\stage_gen[1].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5752_ (.CLK(clknet_3_0__leaf_CLK),
    .D(net501),
    .Q(\stage_gen[1].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5753_ (.CLK(clknet_3_0__leaf_CLK),
    .D(net483),
    .Q(\stage_gen[1].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5754_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net488),
    .Q(\stage_gen[1].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _5755_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_1301_),
    .Q(\stage_gen[1].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _5756_ (.D(_0000_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5757_ (.D(_0001_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5758_ (.D(_0002_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5759_ (.D(_0003_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5760_ (.D(_0004_),
    .GATE_N(net281),
    .Q(\stage_gen[1].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5761_ (.D(_0197_),
    .GATE_N(net368),
    .Q(\stage_gen[1].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5762_ (.D(_0198_),
    .GATE_N(net277),
    .Q(\stage_gen[1].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5763_ (.D(_0199_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5764_ (.D(_0200_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5765_ (.D(_0201_),
    .GATE_N(net282),
    .Q(\stage_gen[1].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5766_ (.D(_0252_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5767_ (.D(_0253_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5768_ (.D(_0254_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5769_ (.D(_0255_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5770_ (.D(_0256_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5771_ (.D(_0307_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5772_ (.D(_0308_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5773_ (.D(_0309_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5774_ (.D(_0310_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5775_ (.D(_0311_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5776_ (.D(_0362_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[4].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5777_ (.D(_0363_),
    .GATE_N(net277),
    .Q(\stage_gen[1].mux_gen[4].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5778_ (.D(_0364_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[4].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5779_ (.D(_0365_),
    .GATE_N(net368),
    .Q(\stage_gen[1].mux_gen[4].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5780_ (.D(_0366_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[4].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5781_ (.D(_0417_),
    .GATE_N(net361),
    .Q(\stage_gen[1].mux_gen[5].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5782_ (.D(_0418_),
    .GATE_N(net277),
    .Q(\stage_gen[1].mux_gen[5].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5783_ (.D(_0419_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[5].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5784_ (.D(_0420_),
    .GATE_N(net368),
    .Q(\stage_gen[1].mux_gen[5].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5785_ (.D(_0421_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[5].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5786_ (.D(_0472_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[6].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5787_ (.D(_0473_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[6].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5788_ (.D(_0474_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[6].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5789_ (.D(_0475_),
    .GATE_N(net361),
    .Q(\stage_gen[1].mux_gen[6].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5790_ (.D(_0476_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[6].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5791_ (.D(_0527_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[7].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5792_ (.D(_0528_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[7].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5793_ (.D(_0529_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[7].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5794_ (.D(_0530_),
    .GATE_N(net361),
    .Q(\stage_gen[1].mux_gen[7].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5795_ (.D(_0531_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[7].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5796_ (.D(_0582_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[8].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5797_ (.D(_0583_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[8].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5798_ (.D(_0584_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[8].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5799_ (.D(_0585_),
    .GATE_N(net361),
    .Q(\stage_gen[1].mux_gen[8].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5800_ (.D(_0586_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[8].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5801_ (.D(_0637_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[9].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5802_ (.D(_0638_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[9].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5803_ (.D(_0639_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[9].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5804_ (.D(_0640_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[9].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5805_ (.D(_0641_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[9].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5806_ (.D(_0057_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[10].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5807_ (.D(_0058_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[10].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5808_ (.D(_0059_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[10].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5809_ (.D(_0060_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[10].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5810_ (.D(_0061_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[10].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5811_ (.D(_0112_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[11].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5812_ (.D(_0113_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[11].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5813_ (.D(_0114_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[11].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5814_ (.D(_0115_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[11].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5815_ (.D(_0116_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[11].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5816_ (.D(_0157_),
    .GATE_N(net336),
    .Q(\stage_gen[1].mux_gen[12].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5817_ (.D(_0158_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[12].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5818_ (.D(_0159_),
    .GATE_N(net336),
    .Q(\stage_gen[1].mux_gen[12].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5819_ (.D(_0160_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[12].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5820_ (.D(_0161_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[12].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5821_ (.D(_0162_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[13].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5822_ (.D(_0163_),
    .GATE_N(net264),
    .Q(\stage_gen[1].mux_gen[13].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5823_ (.D(_0164_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[13].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5824_ (.D(_0165_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[13].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5825_ (.D(_0166_),
    .GATE_N(net264),
    .Q(\stage_gen[1].mux_gen[13].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5826_ (.D(_0167_),
    .GATE_N(net336),
    .Q(\stage_gen[1].mux_gen[14].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5827_ (.D(_0168_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[14].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5828_ (.D(_0169_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[14].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5829_ (.D(_0170_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[14].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5830_ (.D(_0171_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[14].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5831_ (.D(_0172_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[15].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5832_ (.D(_0173_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[15].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5833_ (.D(_0174_),
    .GATE_N(net336),
    .Q(\stage_gen[1].mux_gen[15].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5834_ (.D(_0175_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[15].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5835_ (.D(_0176_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[15].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5836_ (.D(_0177_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[16].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5837_ (.D(_0178_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[16].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5838_ (.D(_0179_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[16].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5839_ (.D(_0180_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[16].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5840_ (.D(_0181_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[16].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5841_ (.D(_0182_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[17].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5842_ (.D(_0183_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[17].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5843_ (.D(_0184_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[17].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5844_ (.D(_0185_),
    .GATE_N(net335),
    .Q(\stage_gen[1].mux_gen[17].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5845_ (.D(_0186_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[17].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5846_ (.D(_0187_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[18].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5847_ (.D(_0188_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[18].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5848_ (.D(_0189_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[18].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5849_ (.D(_0190_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[18].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5850_ (.D(_0191_),
    .GATE_N(net262),
    .Q(\stage_gen[1].mux_gen[18].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5851_ (.D(_0192_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[19].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5852_ (.D(_0193_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[19].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5853_ (.D(_0194_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[19].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5854_ (.D(_0195_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[19].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5855_ (.D(_0196_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[19].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5856_ (.D(_0202_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[20].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5857_ (.D(_0203_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[20].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5858_ (.D(_0204_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[20].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5859_ (.D(_0205_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[20].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5860_ (.D(_0206_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[20].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5861_ (.D(_0207_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[21].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5862_ (.D(_0208_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[21].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5863_ (.D(_0209_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[21].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5864_ (.D(_0210_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[21].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5865_ (.D(_0211_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[21].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5866_ (.D(_0212_),
    .GATE_N(net338),
    .Q(\stage_gen[1].mux_gen[22].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5867_ (.D(_0213_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[22].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5868_ (.D(_0214_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[22].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5869_ (.D(_0215_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[22].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5870_ (.D(_0216_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[22].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5871_ (.D(_0217_),
    .GATE_N(net338),
    .Q(\stage_gen[1].mux_gen[23].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5872_ (.D(_0218_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[23].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5873_ (.D(_0219_),
    .GATE_N(net333),
    .Q(\stage_gen[1].mux_gen[23].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5874_ (.D(_0220_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[23].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5875_ (.D(_0221_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[23].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5876_ (.D(_0222_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[24].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5877_ (.D(_0223_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[24].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5878_ (.D(_0224_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[24].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5879_ (.D(_0225_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[24].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5880_ (.D(_0226_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[24].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5881_ (.D(_0227_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[25].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5882_ (.D(_0228_),
    .GATE_N(net263),
    .Q(\stage_gen[1].mux_gen[25].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5883_ (.D(_0229_),
    .GATE_N(net326),
    .Q(\stage_gen[1].mux_gen[25].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5884_ (.D(_0230_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[25].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5885_ (.D(_0231_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[25].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5886_ (.D(_0232_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[26].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5887_ (.D(_0233_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[26].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5888_ (.D(_0234_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[26].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5889_ (.D(_0235_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[26].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5890_ (.D(_0236_),
    .GATE_N(net261),
    .Q(\stage_gen[1].mux_gen[26].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5891_ (.D(_0237_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[27].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5892_ (.D(_0238_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[27].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5893_ (.D(_0239_),
    .GATE_N(net326),
    .Q(\stage_gen[1].mux_gen[27].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5894_ (.D(_0240_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[27].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5895_ (.D(_0241_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[27].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5896_ (.D(_0242_),
    .GATE_N(net326),
    .Q(\stage_gen[1].mux_gen[28].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5897_ (.D(_0243_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[28].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5898_ (.D(_0244_),
    .GATE_N(net326),
    .Q(\stage_gen[1].mux_gen[28].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5899_ (.D(_0245_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[28].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5900_ (.D(_0246_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[28].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5901_ (.D(_0247_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[29].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5902_ (.D(_0248_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[29].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5903_ (.D(_0249_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[29].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5904_ (.D(_0250_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[29].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5905_ (.D(_0251_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[29].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5906_ (.D(_0257_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[30].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5907_ (.D(_0258_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[30].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5908_ (.D(_0259_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[30].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5909_ (.D(_0260_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[30].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5910_ (.D(_0261_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[30].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5911_ (.D(_0262_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[31].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5912_ (.D(_0263_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[31].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5913_ (.D(_0264_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[31].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5914_ (.D(_0265_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[31].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5915_ (.D(_0266_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[31].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5916_ (.D(_0267_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[32].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5917_ (.D(_0268_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[32].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5918_ (.D(_0269_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[32].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5919_ (.D(_0270_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[32].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5920_ (.D(_0271_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[32].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5921_ (.D(_0272_),
    .GATE_N(net326),
    .Q(\stage_gen[1].mux_gen[33].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5922_ (.D(_0273_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[33].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5923_ (.D(_0274_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[33].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5924_ (.D(_0275_),
    .GATE_N(net325),
    .Q(\stage_gen[1].mux_gen[33].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5925_ (.D(_0276_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[33].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5926_ (.D(_0277_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[34].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5927_ (.D(_0278_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[34].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5928_ (.D(_0279_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[34].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5929_ (.D(_0280_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[34].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5930_ (.D(_0281_),
    .GATE_N(net264),
    .Q(\stage_gen[1].mux_gen[34].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5931_ (.D(_0282_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[35].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5932_ (.D(_0283_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[35].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5933_ (.D(_0284_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[35].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5934_ (.D(_0285_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[35].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5935_ (.D(_0286_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[35].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5936_ (.D(_0287_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[36].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5937_ (.D(_0288_),
    .GATE_N(net259),
    .Q(\stage_gen[1].mux_gen[36].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5938_ (.D(_0289_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[36].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5939_ (.D(_0290_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[36].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5940_ (.D(_0291_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[36].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5941_ (.D(_0292_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[37].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5942_ (.D(_0293_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[37].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5943_ (.D(_0294_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[37].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5944_ (.D(_0295_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[37].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5945_ (.D(_0296_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[37].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5946_ (.D(_0297_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[38].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5947_ (.D(_0298_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[38].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5948_ (.D(_0299_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[38].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5949_ (.D(_0300_),
    .GATE_N(net323),
    .Q(\stage_gen[1].mux_gen[38].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5950_ (.D(_0301_),
    .GATE_N(net260),
    .Q(\stage_gen[1].mux_gen[38].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5951_ (.D(_0302_),
    .GATE_N(net324),
    .Q(\stage_gen[1].mux_gen[39].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5952_ (.D(_0303_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[39].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5953_ (.D(_0304_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[39].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5954_ (.D(_0305_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[39].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5955_ (.D(_0306_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[39].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5956_ (.D(_0312_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[40].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5957_ (.D(_0313_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[40].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5958_ (.D(_0314_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[40].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5959_ (.D(_0315_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[40].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5960_ (.D(_0316_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[40].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5961_ (.D(_0317_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[41].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5962_ (.D(_0318_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[41].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5963_ (.D(_0319_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[41].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5964_ (.D(_0320_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[41].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5965_ (.D(_0321_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[41].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5966_ (.D(_0322_),
    .GATE_N(net331),
    .Q(\stage_gen[1].mux_gen[42].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5967_ (.D(_0323_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[42].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5968_ (.D(_0324_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[42].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5969_ (.D(_0325_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[42].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5970_ (.D(_0326_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[42].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5971_ (.D(_0327_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[43].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5972_ (.D(_0328_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[43].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5973_ (.D(_0329_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[43].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5974_ (.D(_0330_),
    .GATE_N(net331),
    .Q(\stage_gen[1].mux_gen[43].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5975_ (.D(_0331_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[43].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5976_ (.D(_0332_),
    .GATE_N(net328),
    .Q(\stage_gen[1].mux_gen[44].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5977_ (.D(_0333_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[44].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5978_ (.D(_0334_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[44].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5979_ (.D(_0335_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[44].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5980_ (.D(_0336_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[44].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5981_ (.D(_0337_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[45].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5982_ (.D(_0338_),
    .GATE_N(net265),
    .Q(\stage_gen[1].mux_gen[45].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5983_ (.D(_0339_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[45].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5984_ (.D(_0340_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[45].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5985_ (.D(_0341_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[45].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5986_ (.D(_0342_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[46].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5987_ (.D(_0343_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[46].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5988_ (.D(_0344_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[46].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5989_ (.D(_0345_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[46].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5990_ (.D(_0346_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[46].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5991_ (.D(_0347_),
    .GATE_N(net331),
    .Q(\stage_gen[1].mux_gen[47].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5992_ (.D(_0348_),
    .GATE_N(net266),
    .Q(\stage_gen[1].mux_gen[47].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5993_ (.D(_0349_),
    .GATE_N(net331),
    .Q(\stage_gen[1].mux_gen[47].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5994_ (.D(_0350_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[47].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _5995_ (.D(_0351_),
    .GATE_N(net267),
    .Q(\stage_gen[1].mux_gen[47].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _5996_ (.D(_0352_),
    .GATE_N(net344),
    .Q(\stage_gen[1].mux_gen[48].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _5997_ (.D(_0353_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[48].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _5998_ (.D(_0354_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[48].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _5999_ (.D(_0355_),
    .GATE_N(net329),
    .Q(\stage_gen[1].mux_gen[48].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6000_ (.D(_0356_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[48].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6001_ (.D(_0357_),
    .GATE_N(net344),
    .Q(\stage_gen[1].mux_gen[49].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6002_ (.D(_0358_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[49].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6003_ (.D(_0359_),
    .GATE_N(net344),
    .Q(\stage_gen[1].mux_gen[49].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6004_ (.D(_0360_),
    .GATE_N(net344),
    .Q(\stage_gen[1].mux_gen[49].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6005_ (.D(_0361_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[49].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6006_ (.D(_0367_),
    .GATE_N(net327),
    .Q(\stage_gen[1].mux_gen[50].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6007_ (.D(_0368_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[50].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6008_ (.D(_0369_),
    .GATE_N(net346),
    .Q(\stage_gen[1].mux_gen[50].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6009_ (.D(_0370_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[50].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6010_ (.D(_0371_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[50].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6011_ (.D(_0372_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[51].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6012_ (.D(_0373_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[51].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6013_ (.D(_0374_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[51].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6014_ (.D(_0375_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[51].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6015_ (.D(_0376_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[51].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6016_ (.D(_0377_),
    .GATE_N(net346),
    .Q(\stage_gen[1].mux_gen[52].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6017_ (.D(_0378_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[52].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6018_ (.D(_0379_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[52].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6019_ (.D(_0380_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[52].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6020_ (.D(_0381_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[52].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6021_ (.D(_0382_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[53].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6022_ (.D(_0383_),
    .GATE_N(net286),
    .Q(\stage_gen[1].mux_gen[53].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6023_ (.D(_0384_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[53].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6024_ (.D(_0385_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[53].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6025_ (.D(_0386_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[53].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6026_ (.D(_0387_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[54].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6027_ (.D(_0388_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[54].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6028_ (.D(_0389_),
    .GATE_N(net349),
    .Q(\stage_gen[1].mux_gen[54].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6029_ (.D(_0390_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[54].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6030_ (.D(_0391_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[54].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6031_ (.D(_0392_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[55].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6032_ (.D(_0393_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[55].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6033_ (.D(_0394_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[55].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6034_ (.D(_0395_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[55].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6035_ (.D(_0396_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[55].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6036_ (.D(_0397_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[56].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6037_ (.D(_0398_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[56].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6038_ (.D(_0399_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[56].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6039_ (.D(_0400_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[56].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6040_ (.D(_0401_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[56].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6041_ (.D(_0402_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[57].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6042_ (.D(_0403_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[57].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6043_ (.D(_0404_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[57].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6044_ (.D(_0405_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[57].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6045_ (.D(_0406_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[57].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6046_ (.D(_0407_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[58].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6047_ (.D(_0408_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[58].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6048_ (.D(_0409_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[58].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6049_ (.D(_0410_),
    .GATE_N(net346),
    .Q(\stage_gen[1].mux_gen[58].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6050_ (.D(_0411_),
    .GATE_N(net286),
    .Q(\stage_gen[1].mux_gen[58].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6051_ (.D(_0412_),
    .GATE_N(net349),
    .Q(\stage_gen[1].mux_gen[59].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6052_ (.D(_0413_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[59].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6053_ (.D(_0414_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[59].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6054_ (.D(_0415_),
    .GATE_N(net352),
    .Q(\stage_gen[1].mux_gen[59].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6055_ (.D(_0416_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[59].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6056_ (.D(_0422_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[60].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6057_ (.D(_0423_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[60].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6058_ (.D(_0424_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[60].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6059_ (.D(_0425_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[60].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6060_ (.D(_0426_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[60].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6061_ (.D(_0427_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[61].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6062_ (.D(_0428_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[61].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6063_ (.D(_0429_),
    .GATE_N(net349),
    .Q(\stage_gen[1].mux_gen[61].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6064_ (.D(_0430_),
    .GATE_N(net352),
    .Q(\stage_gen[1].mux_gen[61].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6065_ (.D(_0431_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[61].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6066_ (.D(_0432_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[62].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6067_ (.D(_0433_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[62].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6068_ (.D(_0434_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[62].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6069_ (.D(_0435_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[62].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6070_ (.D(_0436_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[62].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6071_ (.D(_0437_),
    .GATE_N(net344),
    .Q(\stage_gen[1].mux_gen[63].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6072_ (.D(_0438_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[63].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6073_ (.D(_0439_),
    .GATE_N(net349),
    .Q(\stage_gen[1].mux_gen[63].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6074_ (.D(_0440_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[63].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6075_ (.D(_0441_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[63].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6076_ (.D(_0442_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[64].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6077_ (.D(_0443_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[64].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6078_ (.D(_0444_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[64].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6079_ (.D(_0445_),
    .GATE_N(net352),
    .Q(\stage_gen[1].mux_gen[64].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6080_ (.D(_0446_),
    .GATE_N(net292),
    .Q(\stage_gen[1].mux_gen[64].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6081_ (.D(_0447_),
    .GATE_N(net350),
    .Q(\stage_gen[1].mux_gen[65].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6082_ (.D(_0448_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[65].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6083_ (.D(_0449_),
    .GATE_N(net348),
    .Q(\stage_gen[1].mux_gen[65].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6084_ (.D(_0450_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[65].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6085_ (.D(_0451_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[65].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6086_ (.D(_0452_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[66].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6087_ (.D(_0453_),
    .GATE_N(net290),
    .Q(\stage_gen[1].mux_gen[66].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6088_ (.D(_0454_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[66].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6089_ (.D(_0455_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[66].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6090_ (.D(_0456_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[66].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6091_ (.D(_0457_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[67].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6092_ (.D(_0458_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[67].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6093_ (.D(_0459_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[67].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6094_ (.D(_0460_),
    .GATE_N(net343),
    .Q(\stage_gen[1].mux_gen[67].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6095_ (.D(_0461_),
    .GATE_N(net285),
    .Q(\stage_gen[1].mux_gen[67].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6096_ (.D(_0462_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[68].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6097_ (.D(_0463_),
    .GATE_N(net286),
    .Q(\stage_gen[1].mux_gen[68].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6098_ (.D(_0464_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[68].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6099_ (.D(_0465_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[68].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6100_ (.D(_0466_),
    .GATE_N(net289),
    .Q(\stage_gen[1].mux_gen[68].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6101_ (.D(_0467_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[69].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6102_ (.D(_0468_),
    .GATE_N(net286),
    .Q(\stage_gen[1].mux_gen[69].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6103_ (.D(_0469_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[69].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6104_ (.D(_0470_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[69].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6105_ (.D(_0471_),
    .GATE_N(net292),
    .Q(\stage_gen[1].mux_gen[69].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6106_ (.D(_0477_),
    .GATE_N(net345),
    .Q(\stage_gen[1].mux_gen[70].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6107_ (.D(_0478_),
    .GATE_N(net286),
    .Q(\stage_gen[1].mux_gen[70].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6108_ (.D(_0479_),
    .GATE_N(net355),
    .Q(\stage_gen[1].mux_gen[70].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6109_ (.D(_0480_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[70].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6110_ (.D(_0481_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[70].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6111_ (.D(_0482_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[71].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6112_ (.D(_0483_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[71].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6113_ (.D(_0484_),
    .GATE_N(net355),
    .Q(\stage_gen[1].mux_gen[71].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6114_ (.D(_0485_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[71].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6115_ (.D(_0486_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[71].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6116_ (.D(_0487_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[72].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6117_ (.D(_0488_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[72].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6118_ (.D(_0489_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[72].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6119_ (.D(_0490_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[72].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6120_ (.D(_0491_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[72].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6121_ (.D(_0492_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[73].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6122_ (.D(_0493_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[73].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6123_ (.D(_0494_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[73].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6124_ (.D(_0495_),
    .GATE_N(net351),
    .Q(\stage_gen[1].mux_gen[73].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6125_ (.D(_0496_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[73].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6126_ (.D(_0497_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[74].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6127_ (.D(_0498_),
    .GATE_N(net284),
    .Q(\stage_gen[1].mux_gen[74].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6128_ (.D(_0499_),
    .GATE_N(net358),
    .Q(\stage_gen[1].mux_gen[74].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6129_ (.D(_0500_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[74].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6130_ (.D(_0501_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[74].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6131_ (.D(_0502_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[75].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6132_ (.D(_0503_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[75].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6133_ (.D(_0504_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[75].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6134_ (.D(_0505_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[75].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6135_ (.D(_0506_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[75].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6136_ (.D(_0507_),
    .GATE_N(net347),
    .Q(\stage_gen[1].mux_gen[76].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6137_ (.D(_0508_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[76].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6138_ (.D(_0509_),
    .GATE_N(net355),
    .Q(\stage_gen[1].mux_gen[76].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6139_ (.D(_0510_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[76].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6140_ (.D(_0511_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[76].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6141_ (.D(_0512_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[77].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6142_ (.D(_0513_),
    .GATE_N(net288),
    .Q(\stage_gen[1].mux_gen[77].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6143_ (.D(_0514_),
    .GATE_N(net355),
    .Q(\stage_gen[1].mux_gen[77].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6144_ (.D(_0515_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[77].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6145_ (.D(_0516_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[77].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6146_ (.D(_0517_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[78].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6147_ (.D(_0518_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[78].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6148_ (.D(_0519_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[78].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6149_ (.D(_0520_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[78].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6150_ (.D(_0521_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[78].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6151_ (.D(_0522_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[79].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6152_ (.D(_0523_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[79].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6153_ (.D(_0524_),
    .GATE_N(net355),
    .Q(\stage_gen[1].mux_gen[79].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6154_ (.D(_0525_),
    .GATE_N(net358),
    .Q(\stage_gen[1].mux_gen[79].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6155_ (.D(_0526_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[79].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6156_ (.D(_0532_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[80].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6157_ (.D(_0533_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[80].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6158_ (.D(_0534_),
    .GATE_N(net354),
    .Q(\stage_gen[1].mux_gen[80].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6159_ (.D(_0535_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[80].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6160_ (.D(_0536_),
    .GATE_N(net292),
    .Q(\stage_gen[1].mux_gen[80].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6161_ (.D(_0537_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[81].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6162_ (.D(_0538_),
    .GATE_N(net283),
    .Q(\stage_gen[1].mux_gen[81].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6163_ (.D(_0539_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[81].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6164_ (.D(_0540_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[81].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6165_ (.D(_0541_),
    .GATE_N(net271),
    .Q(\stage_gen[1].mux_gen[81].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6166_ (.D(_0542_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[82].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6167_ (.D(_0543_),
    .GATE_N(net283),
    .Q(\stage_gen[1].mux_gen[82].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6168_ (.D(_0544_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[82].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6169_ (.D(_0545_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[82].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6170_ (.D(_0546_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[82].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6171_ (.D(_0547_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[83].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6172_ (.D(_0548_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[83].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6173_ (.D(_0549_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[83].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6174_ (.D(_0550_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[83].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6175_ (.D(_0551_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[83].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6176_ (.D(_0552_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[84].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6177_ (.D(_0553_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[84].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6178_ (.D(_0554_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[84].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6179_ (.D(_0555_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[84].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6180_ (.D(_0556_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[84].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6181_ (.D(_0557_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[85].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6182_ (.D(_0558_),
    .GATE_N(net271),
    .Q(\stage_gen[1].mux_gen[85].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6183_ (.D(_0559_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[85].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6184_ (.D(_0560_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[85].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6185_ (.D(_0561_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[85].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6186_ (.D(_0562_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[86].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6187_ (.D(_0563_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[86].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6188_ (.D(_0564_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[86].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6189_ (.D(_0565_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[86].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6190_ (.D(_0566_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[86].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6191_ (.D(_0567_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[87].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6192_ (.D(_0568_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[87].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6193_ (.D(_0569_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[87].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6194_ (.D(_0570_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[87].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6195_ (.D(_0571_),
    .GATE_N(net293),
    .Q(\stage_gen[1].mux_gen[87].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6196_ (.D(_0572_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[88].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6197_ (.D(_0573_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[88].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6198_ (.D(_0574_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[88].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6199_ (.D(_0575_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[88].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6200_ (.D(_0576_),
    .GATE_N(net271),
    .Q(\stage_gen[1].mux_gen[88].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6201_ (.D(_0577_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[89].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6202_ (.D(_0578_),
    .GATE_N(net271),
    .Q(\stage_gen[1].mux_gen[89].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6203_ (.D(_0579_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[89].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6204_ (.D(_0580_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[89].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6205_ (.D(_0581_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[89].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6206_ (.D(_0587_),
    .GATE_N(net375),
    .Q(\stage_gen[1].mux_gen[90].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6207_ (.D(_0588_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[90].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6208_ (.D(_0589_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[90].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6209_ (.D(_0590_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[90].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6210_ (.D(_0591_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[90].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6211_ (.D(_0592_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[91].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6212_ (.D(_0593_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[91].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6213_ (.D(_0594_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[91].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6214_ (.D(_0595_),
    .GATE_N(net330),
    .Q(\stage_gen[1].mux_gen[91].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6215_ (.D(_0596_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[91].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6216_ (.D(_0597_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[92].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6217_ (.D(_0598_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[92].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6218_ (.D(_0599_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[92].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6219_ (.D(_0600_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[92].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6220_ (.D(_0601_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[92].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6221_ (.D(_0602_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[93].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6222_ (.D(_0603_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[93].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6223_ (.D(_0604_),
    .GATE_N(net356),
    .Q(\stage_gen[1].mux_gen[93].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6224_ (.D(_0605_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[93].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6225_ (.D(_0606_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[93].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6226_ (.D(_0607_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[94].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6227_ (.D(_0608_),
    .GATE_N(net287),
    .Q(\stage_gen[1].mux_gen[94].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6228_ (.D(_0609_),
    .GATE_N(net353),
    .Q(\stage_gen[1].mux_gen[94].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6229_ (.D(_0610_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[94].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6230_ (.D(_0611_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[94].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6231_ (.D(_0612_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[95].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6232_ (.D(_0613_),
    .GATE_N(net271),
    .Q(\stage_gen[1].mux_gen[95].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6233_ (.D(_0614_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[95].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6234_ (.D(_0615_),
    .GATE_N(net357),
    .Q(\stage_gen[1].mux_gen[95].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6235_ (.D(_0616_),
    .GATE_N(net291),
    .Q(\stage_gen[1].mux_gen[95].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6236_ (.D(_0617_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[96].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6237_ (.D(_0618_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[96].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6238_ (.D(_0619_),
    .GATE_N(net338),
    .Q(\stage_gen[1].mux_gen[96].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6239_ (.D(_0620_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[96].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6240_ (.D(_0621_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[96].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6241_ (.D(_0622_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[97].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6242_ (.D(_0623_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[97].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6243_ (.D(_0624_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[97].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6244_ (.D(_0625_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[97].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6245_ (.D(_0626_),
    .GATE_N(net269),
    .Q(\stage_gen[1].mux_gen[97].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6246_ (.D(_0627_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[98].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6247_ (.D(_0628_),
    .GATE_N(net270),
    .Q(\stage_gen[1].mux_gen[98].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6248_ (.D(_0629_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[98].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6249_ (.D(_0630_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[98].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6250_ (.D(_0631_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[98].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6251_ (.D(_0632_),
    .GATE_N(net340),
    .Q(\stage_gen[1].mux_gen[99].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6252_ (.D(_0633_),
    .GATE_N(net269),
    .Q(\stage_gen[1].mux_gen[99].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6253_ (.D(_0634_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[99].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6254_ (.D(_0635_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[99].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6255_ (.D(_0636_),
    .GATE_N(net282),
    .Q(\stage_gen[1].mux_gen[99].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6256_ (.D(_0007_),
    .GATE_N(net339),
    .Q(\stage_gen[1].mux_gen[100].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6257_ (.D(_0008_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[100].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6258_ (.D(_0009_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[100].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6259_ (.D(_0010_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[100].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6260_ (.D(_0011_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[100].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6261_ (.D(_0012_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[101].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6262_ (.D(_0013_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[101].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6263_ (.D(_0014_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[101].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6264_ (.D(_0015_),
    .GATE_N(net338),
    .Q(\stage_gen[1].mux_gen[101].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6265_ (.D(_0016_),
    .GATE_N(net269),
    .Q(\stage_gen[1].mux_gen[101].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6266_ (.D(_0017_),
    .GATE_N(net334),
    .Q(\stage_gen[1].mux_gen[102].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6267_ (.D(_0018_),
    .GATE_N(net269),
    .Q(\stage_gen[1].mux_gen[102].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6268_ (.D(_0019_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[102].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6269_ (.D(_0020_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[102].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6270_ (.D(_0021_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[102].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6271_ (.D(_0022_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[103].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6272_ (.D(_0023_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[103].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6273_ (.D(_0024_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[103].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6274_ (.D(_0025_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[103].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6275_ (.D(_0026_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[103].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6276_ (.D(_0027_),
    .GATE_N(net338),
    .Q(\stage_gen[1].mux_gen[104].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6277_ (.D(_0028_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[104].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6278_ (.D(_0029_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[104].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6279_ (.D(_0030_),
    .GATE_N(net337),
    .Q(\stage_gen[1].mux_gen[104].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6280_ (.D(_0031_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[104].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6281_ (.D(_0032_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[105].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6282_ (.D(_0033_),
    .GATE_N(net283),
    .Q(\stage_gen[1].mux_gen[105].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6283_ (.D(_0034_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[105].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6284_ (.D(_0035_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[105].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6285_ (.D(_0036_),
    .GATE_N(net282),
    .Q(\stage_gen[1].mux_gen[105].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6286_ (.D(_0037_),
    .GATE_N(net332),
    .Q(\stage_gen[1].mux_gen[106].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6287_ (.D(_0038_),
    .GATE_N(net268),
    .Q(\stage_gen[1].mux_gen[106].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6288_ (.D(_0039_),
    .GATE_N(net341),
    .Q(\stage_gen[1].mux_gen[106].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6289_ (.D(_0040_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[106].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6290_ (.D(_0041_),
    .GATE_N(net269),
    .Q(\stage_gen[1].mux_gen[106].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6291_ (.D(_0042_),
    .GATE_N(net365),
    .Q(\stage_gen[1].mux_gen[107].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6292_ (.D(_0043_),
    .GATE_N(net283),
    .Q(\stage_gen[1].mux_gen[107].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6293_ (.D(_0044_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[107].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6294_ (.D(_0045_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[107].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6295_ (.D(_0046_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[107].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6296_ (.D(_0047_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[108].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6297_ (.D(_0048_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[108].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6298_ (.D(_0049_),
    .GATE_N(net374),
    .Q(\stage_gen[1].mux_gen[108].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6299_ (.D(_0050_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[108].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6300_ (.D(_0051_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[108].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6301_ (.D(_0052_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[109].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6302_ (.D(_0053_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[109].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6303_ (.D(_0054_),
    .GATE_N(net370),
    .Q(\stage_gen[1].mux_gen[109].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6304_ (.D(_0055_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[109].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6305_ (.D(_0056_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[109].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6306_ (.D(_0062_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[110].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6307_ (.D(_0063_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[110].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6308_ (.D(_0064_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[110].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6309_ (.D(_0065_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[110].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6310_ (.D(_0066_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[110].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6311_ (.D(_0067_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[111].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6312_ (.D(_0068_),
    .GATE_N(net281),
    .Q(\stage_gen[1].mux_gen[111].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6313_ (.D(_0069_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[111].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6314_ (.D(_0070_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[111].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6315_ (.D(_0071_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[111].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6316_ (.D(_0072_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[112].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6317_ (.D(_0073_),
    .GATE_N(net278),
    .Q(\stage_gen[1].mux_gen[112].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6318_ (.D(_0074_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[112].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6319_ (.D(_0075_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[112].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6320_ (.D(_0076_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[112].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6321_ (.D(_0077_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[113].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6322_ (.D(_0078_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[113].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6323_ (.D(_0079_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[113].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6324_ (.D(_0080_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[113].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6325_ (.D(_0081_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[113].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6326_ (.D(_0082_),
    .GATE_N(net367),
    .Q(\stage_gen[1].mux_gen[114].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6327_ (.D(_0083_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[114].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6328_ (.D(_0084_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[114].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6329_ (.D(_0085_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[114].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6330_ (.D(_0086_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[114].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6331_ (.D(_0087_),
    .GATE_N(net362),
    .Q(\stage_gen[1].mux_gen[115].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6332_ (.D(_0088_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[115].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6333_ (.D(_0089_),
    .GATE_N(net362),
    .Q(\stage_gen[1].mux_gen[115].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6334_ (.D(_0090_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[115].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6335_ (.D(_0091_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[115].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6336_ (.D(_0092_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[116].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6337_ (.D(_0093_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[116].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6338_ (.D(_0094_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[116].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6339_ (.D(_0095_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[116].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6340_ (.D(_0096_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[116].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6341_ (.D(_0097_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[117].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6342_ (.D(_0098_),
    .GATE_N(net281),
    .Q(\stage_gen[1].mux_gen[117].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6343_ (.D(_0099_),
    .GATE_N(net373),
    .Q(\stage_gen[1].mux_gen[117].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6344_ (.D(_0100_),
    .GATE_N(net374),
    .Q(\stage_gen[1].mux_gen[117].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6345_ (.D(_0101_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[117].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6346_ (.D(_0102_),
    .GATE_N(net368),
    .Q(\stage_gen[1].mux_gen[118].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6347_ (.D(_0103_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[118].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6348_ (.D(_0104_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[118].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6349_ (.D(_0105_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[118].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6350_ (.D(_0106_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[118].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6351_ (.D(_0107_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[119].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6352_ (.D(_0108_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[119].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6353_ (.D(_0109_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[119].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6354_ (.D(_0110_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[119].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6355_ (.D(_0111_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[119].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6356_ (.D(_0117_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[120].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6357_ (.D(_0118_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[120].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6358_ (.D(_0119_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[120].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6359_ (.D(_0120_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[120].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6360_ (.D(_0121_),
    .GATE_N(net279),
    .Q(\stage_gen[1].mux_gen[120].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6361_ (.D(_0122_),
    .GATE_N(net336),
    .Q(\stage_gen[1].mux_gen[121].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6362_ (.D(_0123_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[121].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6363_ (.D(_0124_),
    .GATE_N(net362),
    .Q(\stage_gen[1].mux_gen[121].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6364_ (.D(_0125_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[121].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6365_ (.D(_0126_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[121].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6366_ (.D(_0127_),
    .GATE_N(net371),
    .Q(\stage_gen[1].mux_gen[122].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6367_ (.D(_0128_),
    .GATE_N(net280),
    .Q(\stage_gen[1].mux_gen[122].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6368_ (.D(_0129_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[122].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6369_ (.D(_0130_),
    .GATE_N(net372),
    .Q(\stage_gen[1].mux_gen[122].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6370_ (.D(_0131_),
    .GATE_N(net281),
    .Q(\stage_gen[1].mux_gen[122].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6371_ (.D(_0132_),
    .GATE_N(net361),
    .Q(\stage_gen[1].mux_gen[123].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6372_ (.D(_0133_),
    .GATE_N(net277),
    .Q(\stage_gen[1].mux_gen[123].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6373_ (.D(_0134_),
    .GATE_N(net370),
    .Q(\stage_gen[1].mux_gen[123].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6374_ (.D(_0135_),
    .GATE_N(net368),
    .Q(\stage_gen[1].mux_gen[123].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6375_ (.D(_0136_),
    .GATE_N(net276),
    .Q(\stage_gen[1].mux_gen[123].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6376_ (.D(_0137_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[124].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6377_ (.D(_0138_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[124].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6378_ (.D(_0139_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[124].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6379_ (.D(_0140_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[124].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6380_ (.D(_0141_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[124].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6381_ (.D(_0142_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[125].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6382_ (.D(_0143_),
    .GATE_N(net273),
    .Q(\stage_gen[1].mux_gen[125].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6383_ (.D(_0144_),
    .GATE_N(net360),
    .Q(\stage_gen[1].mux_gen[125].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6384_ (.D(_0145_),
    .GATE_N(net363),
    .Q(\stage_gen[1].mux_gen[125].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6385_ (.D(_0146_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[125].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6386_ (.D(_0147_),
    .GATE_N(net366),
    .Q(\stage_gen[1].mux_gen[126].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6387_ (.D(_0148_),
    .GATE_N(net275),
    .Q(\stage_gen[1].mux_gen[126].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6388_ (.D(_0149_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[126].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6389_ (.D(_0150_),
    .GATE_N(net369),
    .Q(\stage_gen[1].mux_gen[126].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6390_ (.D(_0151_),
    .GATE_N(net278),
    .Q(\stage_gen[1].mux_gen[126].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6391_ (.D(_0152_),
    .GATE_N(net364),
    .Q(\stage_gen[1].mux_gen[127].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6392_ (.D(_0153_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[127].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6393_ (.D(_0154_),
    .GATE_N(net362),
    .Q(\stage_gen[1].mux_gen[127].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6394_ (.D(_0155_),
    .GATE_N(net359),
    .Q(\stage_gen[1].mux_gen[127].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6395_ (.D(_0156_),
    .GATE_N(net274),
    .Q(\stage_gen[1].mux_gen[127].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _6396_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_1302_),
    .Q(\stage_gen[2].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6397_ (.CLK(clknet_3_4__leaf_CLK),
    .D(net511),
    .Q(\stage_gen[2].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6398_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net512),
    .Q(\stage_gen[2].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6399_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_1305_),
    .Q(\stage_gen[2].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6400_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net517),
    .Q(\stage_gen[2].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6401_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net502),
    .Q(\stage_gen[2].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6402_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net489),
    .Q(\stage_gen[2].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6403_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net503),
    .Q(\stage_gen[2].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6404_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net490),
    .Q(\stage_gen[2].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6405_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net491),
    .Q(\stage_gen[2].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6406_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_1312_),
    .Q(\stage_gen[2].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _6407_ (.D(_0642_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6408_ (.D(_0643_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6409_ (.D(_0644_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6410_ (.D(_0645_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6411_ (.D(_0646_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6412_ (.D(_0699_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6413_ (.D(_0700_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6414_ (.D(_0701_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6415_ (.D(_0702_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6416_ (.D(_0703_),
    .GATE_N(net311),
    .Q(\stage_gen[2].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6417_ (.D(_0754_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6418_ (.D(_0755_),
    .GATE_N(net311),
    .Q(\stage_gen[2].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6419_ (.D(_0756_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6420_ (.D(_0757_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6421_ (.D(_0758_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6422_ (.D(_0809_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6423_ (.D(_0810_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6424_ (.D(_0811_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6425_ (.D(_0812_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6426_ (.D(_0813_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6427_ (.D(_0864_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[4].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6428_ (.D(_0865_),
    .GATE_N(net309),
    .Q(\stage_gen[2].mux_gen[4].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6429_ (.D(_0866_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[4].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6430_ (.D(_0867_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[4].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6431_ (.D(_0868_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[4].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6432_ (.D(_0919_),
    .GATE_N(net411),
    .Q(\stage_gen[2].mux_gen[5].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6433_ (.D(_0920_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[5].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6434_ (.D(_0921_),
    .GATE_N(net411),
    .Q(\stage_gen[2].mux_gen[5].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6435_ (.D(_0922_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[5].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6436_ (.D(_0923_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[5].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6437_ (.D(_0944_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[6].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6438_ (.D(_0945_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[6].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6439_ (.D(_0946_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[6].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6440_ (.D(_0947_),
    .GATE_N(net419),
    .Q(\stage_gen[2].mux_gen[6].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6441_ (.D(_0948_),
    .GATE_N(net309),
    .Q(\stage_gen[2].mux_gen[6].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6442_ (.D(_0949_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[7].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6443_ (.D(_0950_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[7].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6444_ (.D(_0951_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[7].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6445_ (.D(_0952_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[7].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6446_ (.D(_0953_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[7].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6447_ (.D(_0954_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[8].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6448_ (.D(_0955_),
    .GATE_N(net309),
    .Q(\stage_gen[2].mux_gen[8].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6449_ (.D(_0956_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[8].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6450_ (.D(_0957_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[8].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6451_ (.D(_0958_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[8].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6452_ (.D(_0959_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[9].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6453_ (.D(_0960_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[9].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6454_ (.D(_0961_),
    .GATE_N(net410),
    .Q(\stage_gen[2].mux_gen[9].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6455_ (.D(_0962_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[9].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6456_ (.D(_0963_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[9].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6457_ (.D(_0649_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[10].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6458_ (.D(_0650_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[10].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6459_ (.D(_0651_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[10].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6460_ (.D(_0652_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[10].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6461_ (.D(_0653_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[10].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6462_ (.D(_0654_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[11].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6463_ (.D(_0655_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[11].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6464_ (.D(_0656_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[11].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6465_ (.D(_0657_),
    .GATE_N(net406),
    .Q(\stage_gen[2].mux_gen[11].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6466_ (.D(_0658_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[11].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6467_ (.D(_0659_),
    .GATE_N(net405),
    .Q(\stage_gen[2].mux_gen[12].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6468_ (.D(_0660_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[12].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6469_ (.D(_0661_),
    .GATE_N(net406),
    .Q(\stage_gen[2].mux_gen[12].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6470_ (.D(_0662_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[12].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6471_ (.D(_0663_),
    .GATE_N(net305),
    .Q(\stage_gen[2].mux_gen[12].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6472_ (.D(_0664_),
    .GATE_N(net404),
    .Q(\stage_gen[2].mux_gen[13].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6473_ (.D(_0665_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[13].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6474_ (.D(_0666_),
    .GATE_N(net404),
    .Q(\stage_gen[2].mux_gen[13].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6475_ (.D(_0667_),
    .GATE_N(net404),
    .Q(\stage_gen[2].mux_gen[13].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6476_ (.D(_0668_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[13].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6477_ (.D(_0669_),
    .GATE_N(net404),
    .Q(\stage_gen[2].mux_gen[14].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6478_ (.D(_0670_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[14].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6479_ (.D(_0671_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[14].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6480_ (.D(_0672_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[14].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6481_ (.D(_0673_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[14].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6482_ (.D(_0674_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[15].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6483_ (.D(_0675_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[15].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6484_ (.D(_0676_),
    .GATE_N(net404),
    .Q(\stage_gen[2].mux_gen[15].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6485_ (.D(_0677_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[15].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6486_ (.D(_0678_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[15].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6487_ (.D(_0679_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[16].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6488_ (.D(_0680_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[16].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6489_ (.D(_0681_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[16].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6490_ (.D(_0682_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[16].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6491_ (.D(_0683_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[16].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6492_ (.D(_0684_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[17].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6493_ (.D(_0685_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[17].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6494_ (.D(_0686_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[17].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6495_ (.D(_0687_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[17].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6496_ (.D(_0688_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[17].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6497_ (.D(_0689_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[18].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6498_ (.D(_0690_),
    .GATE_N(net304),
    .Q(\stage_gen[2].mux_gen[18].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6499_ (.D(_0691_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[18].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6500_ (.D(_0692_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[18].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6501_ (.D(_0693_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[18].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6502_ (.D(_0694_),
    .GATE_N(net403),
    .Q(\stage_gen[2].mux_gen[19].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6503_ (.D(_0695_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[19].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6504_ (.D(_0696_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[19].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6505_ (.D(_0697_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[19].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6506_ (.D(_0698_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[19].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6507_ (.D(_0704_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[20].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6508_ (.D(_0705_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[20].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6509_ (.D(_0706_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[20].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6510_ (.D(_0707_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[20].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6511_ (.D(_0708_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[20].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6512_ (.D(_0709_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[21].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6513_ (.D(_0710_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[21].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6514_ (.D(_0711_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[21].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6515_ (.D(_0712_),
    .GATE_N(net407),
    .Q(\stage_gen[2].mux_gen[21].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6516_ (.D(_0713_),
    .GATE_N(net306),
    .Q(\stage_gen[2].mux_gen[21].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6517_ (.D(_0714_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[22].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6518_ (.D(_0715_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[22].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6519_ (.D(_0716_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[22].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6520_ (.D(_0717_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[22].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6521_ (.D(_0718_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[22].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6522_ (.D(_0719_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[23].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6523_ (.D(_0720_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[23].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6524_ (.D(_0721_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[23].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6525_ (.D(_0722_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[23].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6526_ (.D(_0723_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[23].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6527_ (.D(_0724_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[24].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6528_ (.D(_0725_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[24].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6529_ (.D(_0726_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[24].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6530_ (.D(_0727_),
    .GATE_N(net420),
    .Q(\stage_gen[2].mux_gen[24].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6531_ (.D(_0728_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[24].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6532_ (.D(_0729_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[25].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6533_ (.D(_0730_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[25].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6534_ (.D(_0731_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[25].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6535_ (.D(_0732_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[25].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6536_ (.D(_0733_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[25].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6537_ (.D(_0734_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[26].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6538_ (.D(_0735_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[26].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6539_ (.D(_0736_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[26].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6540_ (.D(_0737_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[26].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6541_ (.D(_0738_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[26].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6542_ (.D(_0739_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[27].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6543_ (.D(_0740_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[27].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6544_ (.D(_0741_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[27].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6545_ (.D(_0742_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[27].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6546_ (.D(_0743_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[27].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6547_ (.D(_0744_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[28].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6548_ (.D(_0745_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[28].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6549_ (.D(_0746_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[28].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6550_ (.D(_0747_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[28].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6551_ (.D(_0748_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[28].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6552_ (.D(_0749_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[29].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6553_ (.D(_0750_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[29].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6554_ (.D(_0751_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[29].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6555_ (.D(_0752_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[29].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6556_ (.D(_0753_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[29].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6557_ (.D(_0759_),
    .GATE_N(net423),
    .Q(\stage_gen[2].mux_gen[30].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6558_ (.D(_0760_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[30].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6559_ (.D(_0761_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[30].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6560_ (.D(_0762_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[30].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6561_ (.D(_0763_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[30].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6562_ (.D(_0764_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[31].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6563_ (.D(_0765_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[31].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6564_ (.D(_0766_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[31].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6565_ (.D(_0767_),
    .GATE_N(net424),
    .Q(\stage_gen[2].mux_gen[31].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6566_ (.D(_0768_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[31].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6567_ (.D(_0769_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[32].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6568_ (.D(_0770_),
    .GATE_N(net317),
    .Q(\stage_gen[2].mux_gen[32].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6569_ (.D(_0771_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[32].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6570_ (.D(_0772_),
    .GATE_N(net423),
    .Q(\stage_gen[2].mux_gen[32].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6571_ (.D(_0773_),
    .GATE_N(net318),
    .Q(\stage_gen[2].mux_gen[32].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6572_ (.D(_0774_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[33].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6573_ (.D(_0775_),
    .GATE_N(net318),
    .Q(\stage_gen[2].mux_gen[33].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6574_ (.D(_0776_),
    .GATE_N(net425),
    .Q(\stage_gen[2].mux_gen[33].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6575_ (.D(_0777_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[33].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6576_ (.D(_0778_),
    .GATE_N(net318),
    .Q(\stage_gen[2].mux_gen[33].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6577_ (.D(_0779_),
    .GATE_N(net423),
    .Q(\stage_gen[2].mux_gen[34].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6578_ (.D(_0780_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[34].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6579_ (.D(_0781_),
    .GATE_N(net422),
    .Q(\stage_gen[2].mux_gen[34].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6580_ (.D(_0782_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[34].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6581_ (.D(_0783_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[34].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6582_ (.D(_0784_),
    .GATE_N(net423),
    .Q(\stage_gen[2].mux_gen[35].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6583_ (.D(_0785_),
    .GATE_N(net318),
    .Q(\stage_gen[2].mux_gen[35].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6584_ (.D(_0786_),
    .GATE_N(net428),
    .Q(\stage_gen[2].mux_gen[35].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6585_ (.D(_0787_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[35].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6586_ (.D(_0788_),
    .GATE_N(net318),
    .Q(\stage_gen[2].mux_gen[35].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6587_ (.D(_0789_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[36].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6588_ (.D(_0790_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[36].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6589_ (.D(_0791_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[36].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6590_ (.D(_0792_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[36].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6591_ (.D(_0793_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[36].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6592_ (.D(_0794_),
    .GATE_N(net423),
    .Q(\stage_gen[2].mux_gen[37].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6593_ (.D(_0795_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[37].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6594_ (.D(_0796_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[37].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6595_ (.D(_0797_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[37].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6596_ (.D(_0798_),
    .GATE_N(net319),
    .Q(\stage_gen[2].mux_gen[37].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6597_ (.D(_0799_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[38].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6598_ (.D(_0800_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[38].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6599_ (.D(_0801_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[38].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6600_ (.D(_0802_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[38].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6601_ (.D(_0803_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[38].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6602_ (.D(_0804_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[39].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6603_ (.D(_0805_),
    .GATE_N(net321),
    .Q(\stage_gen[2].mux_gen[39].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6604_ (.D(_0806_),
    .GATE_N(net430),
    .Q(\stage_gen[2].mux_gen[39].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6605_ (.D(_0807_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[39].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6606_ (.D(_0808_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[39].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6607_ (.D(_0814_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[40].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6608_ (.D(_0815_),
    .GATE_N(net321),
    .Q(\stage_gen[2].mux_gen[40].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6609_ (.D(_0816_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[40].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6610_ (.D(_0817_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[40].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6611_ (.D(_0818_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[40].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6612_ (.D(_0819_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[41].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6613_ (.D(_0820_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[41].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6614_ (.D(_0821_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[41].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6615_ (.D(_0822_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[41].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6616_ (.D(_0823_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[41].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6617_ (.D(_0824_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[42].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6618_ (.D(_0825_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[42].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6619_ (.D(_0826_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[42].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6620_ (.D(_0827_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[42].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6621_ (.D(_0828_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[42].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6622_ (.D(_0829_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[43].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6623_ (.D(_0830_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[43].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6624_ (.D(_0831_),
    .GATE_N(net430),
    .Q(\stage_gen[2].mux_gen[43].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6625_ (.D(_0832_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[43].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6626_ (.D(_0833_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[43].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6627_ (.D(_0834_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[44].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6628_ (.D(_0835_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[44].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6629_ (.D(_0836_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[44].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6630_ (.D(_0837_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[44].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6631_ (.D(_0838_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[44].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6632_ (.D(_0839_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[45].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6633_ (.D(_0840_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[45].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6634_ (.D(_0841_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[45].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6635_ (.D(_0842_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[45].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6636_ (.D(_0843_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[45].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6637_ (.D(_0844_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[46].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6638_ (.D(_0845_),
    .GATE_N(net321),
    .Q(\stage_gen[2].mux_gen[46].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6639_ (.D(_0846_),
    .GATE_N(net427),
    .Q(\stage_gen[2].mux_gen[46].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6640_ (.D(_0847_),
    .GATE_N(net426),
    .Q(\stage_gen[2].mux_gen[46].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6641_ (.D(_0848_),
    .GATE_N(net320),
    .Q(\stage_gen[2].mux_gen[46].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6642_ (.D(_0849_),
    .GATE_N(net421),
    .Q(\stage_gen[2].mux_gen[47].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6643_ (.D(_0850_),
    .GATE_N(net316),
    .Q(\stage_gen[2].mux_gen[47].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6644_ (.D(_0851_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[47].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6645_ (.D(_0852_),
    .GATE_N(net429),
    .Q(\stage_gen[2].mux_gen[47].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6646_ (.D(_0853_),
    .GATE_N(net322),
    .Q(\stage_gen[2].mux_gen[47].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6647_ (.D(_0854_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[48].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6648_ (.D(_0855_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[48].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6649_ (.D(_0856_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[48].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6650_ (.D(_0857_),
    .GATE_N(net417),
    .Q(\stage_gen[2].mux_gen[48].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6651_ (.D(_0858_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[48].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6652_ (.D(_0859_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[49].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6653_ (.D(_0860_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[49].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6654_ (.D(_0861_),
    .GATE_N(net417),
    .Q(\stage_gen[2].mux_gen[49].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6655_ (.D(_0862_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[49].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6656_ (.D(_0863_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[49].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6657_ (.D(_0869_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[50].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6658_ (.D(_0870_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[50].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6659_ (.D(_0871_),
    .GATE_N(net409),
    .Q(\stage_gen[2].mux_gen[50].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6660_ (.D(_0872_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[50].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6661_ (.D(_0873_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[50].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6662_ (.D(_0874_),
    .GATE_N(net409),
    .Q(\stage_gen[2].mux_gen[51].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6663_ (.D(_0875_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[51].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6664_ (.D(_0876_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[51].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6665_ (.D(_0877_),
    .GATE_N(net417),
    .Q(\stage_gen[2].mux_gen[51].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6666_ (.D(_0878_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[51].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6667_ (.D(_0879_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[52].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6668_ (.D(_0880_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[52].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6669_ (.D(_0881_),
    .GATE_N(net409),
    .Q(\stage_gen[2].mux_gen[52].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6670_ (.D(_0882_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[52].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6671_ (.D(_0883_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[52].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6672_ (.D(_0884_),
    .GATE_N(net408),
    .Q(\stage_gen[2].mux_gen[53].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6673_ (.D(_0885_),
    .GATE_N(net307),
    .Q(\stage_gen[2].mux_gen[53].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6674_ (.D(_0886_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[53].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6675_ (.D(_0887_),
    .GATE_N(net417),
    .Q(\stage_gen[2].mux_gen[53].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6676_ (.D(_0888_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[53].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6677_ (.D(_0889_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[54].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6678_ (.D(_0890_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[54].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6679_ (.D(_0891_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[54].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6680_ (.D(_0892_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[54].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6681_ (.D(_0893_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[54].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6682_ (.D(_0894_),
    .GATE_N(net411),
    .Q(\stage_gen[2].mux_gen[55].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6683_ (.D(_0895_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[55].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6684_ (.D(_0896_),
    .GATE_N(net417),
    .Q(\stage_gen[2].mux_gen[55].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6685_ (.D(_0897_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[55].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6686_ (.D(_0898_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[55].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6687_ (.D(_0899_),
    .GATE_N(net411),
    .Q(\stage_gen[2].mux_gen[56].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6688_ (.D(_0900_),
    .GATE_N(net308),
    .Q(\stage_gen[2].mux_gen[56].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6689_ (.D(_0901_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[56].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6690_ (.D(_0902_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[56].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6691_ (.D(_0903_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[56].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6692_ (.D(_0904_),
    .GATE_N(net411),
    .Q(\stage_gen[2].mux_gen[57].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6693_ (.D(_0905_),
    .GATE_N(net309),
    .Q(\stage_gen[2].mux_gen[57].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6694_ (.D(_0906_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[57].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6695_ (.D(_0907_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[57].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6696_ (.D(_0908_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[57].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6697_ (.D(_0909_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[58].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6698_ (.D(_0910_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[58].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6699_ (.D(_0911_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[58].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6700_ (.D(_0912_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[58].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6701_ (.D(_0913_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[58].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6702_ (.D(_0914_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[59].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6703_ (.D(_0915_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[59].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6704_ (.D(_0916_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[59].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6705_ (.D(_0917_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[59].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6706_ (.D(_0918_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[59].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6707_ (.D(_0924_),
    .GATE_N(net416),
    .Q(\stage_gen[2].mux_gen[60].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6708_ (.D(_0925_),
    .GATE_N(net312),
    .Q(\stage_gen[2].mux_gen[60].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6709_ (.D(_0926_),
    .GATE_N(net418),
    .Q(\stage_gen[2].mux_gen[60].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6710_ (.D(_0927_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[60].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6711_ (.D(_0928_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[60].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6712_ (.D(_0929_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[61].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6713_ (.D(_0930_),
    .GATE_N(net311),
    .Q(\stage_gen[2].mux_gen[61].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6714_ (.D(_0931_),
    .GATE_N(net414),
    .Q(\stage_gen[2].mux_gen[61].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6715_ (.D(_0932_),
    .GATE_N(net414),
    .Q(\stage_gen[2].mux_gen[61].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6716_ (.D(_0933_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[61].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6717_ (.D(_0934_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[62].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6718_ (.D(_0935_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[62].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6719_ (.D(_0936_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[62].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6720_ (.D(_0937_),
    .GATE_N(net412),
    .Q(\stage_gen[2].mux_gen[62].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6721_ (.D(_0938_),
    .GATE_N(net313),
    .Q(\stage_gen[2].mux_gen[62].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6722_ (.D(_0939_),
    .GATE_N(net415),
    .Q(\stage_gen[2].mux_gen[63].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6723_ (.D(_0940_),
    .GATE_N(net311),
    .Q(\stage_gen[2].mux_gen[63].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6724_ (.D(_0941_),
    .GATE_N(net413),
    .Q(\stage_gen[2].mux_gen[63].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6725_ (.D(_0942_),
    .GATE_N(net414),
    .Q(\stage_gen[2].mux_gen[63].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6726_ (.D(_0943_),
    .GATE_N(net310),
    .Q(\stage_gen[2].mux_gen[63].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _6727_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_1313_),
    .Q(\stage_gen[3].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6728_ (.CLK(clknet_3_4__leaf_CLK),
    .D(net513),
    .Q(\stage_gen[3].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6729_ (.CLK(clknet_3_5__leaf_CLK),
    .D(net518),
    .Q(\stage_gen[3].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6730_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_1316_),
    .Q(\stage_gen[3].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6731_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net492),
    .Q(\stage_gen[3].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6732_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net504),
    .Q(\stage_gen[3].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6733_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net493),
    .Q(\stage_gen[3].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6734_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net505),
    .Q(\stage_gen[3].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6735_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net479),
    .Q(\stage_gen[3].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6736_ (.CLK(clknet_3_4__leaf_CLK),
    .D(net480),
    .Q(\stage_gen[3].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6737_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_1323_),
    .Q(\stage_gen[3].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _6738_ (.D(_0964_),
    .GATE_N(net395),
    .Q(\stage_gen[3].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6739_ (.D(_0965_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6740_ (.D(_0966_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6741_ (.D(_0967_),
    .GATE_N(net395),
    .Q(\stage_gen[3].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6742_ (.D(_0968_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6743_ (.D(_1021_),
    .GATE_N(net395),
    .Q(\stage_gen[3].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6744_ (.D(_1022_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6745_ (.D(_1023_),
    .GATE_N(net395),
    .Q(\stage_gen[3].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6746_ (.D(_1024_),
    .GATE_N(net395),
    .Q(\stage_gen[3].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6747_ (.D(_1025_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6748_ (.D(_1076_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6749_ (.D(_1077_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6750_ (.D(_1078_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6751_ (.D(_1079_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6752_ (.D(_1080_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6753_ (.D(_1091_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6754_ (.D(_1092_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6755_ (.D(_1093_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6756_ (.D(_1094_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6757_ (.D(_1095_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6758_ (.D(_1096_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[4].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6759_ (.D(_1097_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[4].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6760_ (.D(_1098_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[4].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6761_ (.D(_1099_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[4].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6762_ (.D(_1100_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[4].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6763_ (.D(_1101_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[5].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6764_ (.D(_1102_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[5].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6765_ (.D(_1103_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[5].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6766_ (.D(_1104_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[5].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6767_ (.D(_1105_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[5].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6768_ (.D(_1106_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[6].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6769_ (.D(_1107_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[6].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6770_ (.D(_1108_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[6].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6771_ (.D(_1109_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[6].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6772_ (.D(_1110_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[6].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6773_ (.D(_1111_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[7].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6774_ (.D(_1112_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[7].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6775_ (.D(_1113_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[7].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6776_ (.D(_1114_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[7].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6777_ (.D(_1115_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[7].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6778_ (.D(_1116_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[8].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6779_ (.D(_1117_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[8].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6780_ (.D(_1118_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[8].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6781_ (.D(_1119_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[8].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6782_ (.D(_1120_),
    .GATE_N(net303),
    .Q(\stage_gen[3].mux_gen[8].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6783_ (.D(_1121_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[9].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6784_ (.D(_1122_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[9].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6785_ (.D(_1123_),
    .GATE_N(net389),
    .Q(\stage_gen[3].mux_gen[9].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6786_ (.D(_1124_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[9].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6787_ (.D(_1125_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[9].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6788_ (.D(_0971_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[10].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6789_ (.D(_0972_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[10].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6790_ (.D(_0973_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[10].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6791_ (.D(_0974_),
    .GATE_N(net393),
    .Q(\stage_gen[3].mux_gen[10].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6792_ (.D(_0975_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[10].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6793_ (.D(_0976_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[11].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6794_ (.D(_0977_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[11].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6795_ (.D(_0978_),
    .GATE_N(net389),
    .Q(\stage_gen[3].mux_gen[11].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6796_ (.D(_0979_),
    .GATE_N(net389),
    .Q(\stage_gen[3].mux_gen[11].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6797_ (.D(_0980_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[11].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6798_ (.D(_0981_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[12].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6799_ (.D(_0982_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[12].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6800_ (.D(_0983_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[12].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6801_ (.D(_0984_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[12].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6802_ (.D(_0985_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[12].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6803_ (.D(_0986_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[13].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6804_ (.D(_0987_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[13].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6805_ (.D(_0988_),
    .GATE_N(net389),
    .Q(\stage_gen[3].mux_gen[13].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6806_ (.D(_0989_),
    .GATE_N(net393),
    .Q(\stage_gen[3].mux_gen[13].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6807_ (.D(_0990_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[13].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6808_ (.D(_0991_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[14].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6809_ (.D(_0992_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[14].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6810_ (.D(_0993_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[14].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6811_ (.D(_0994_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[14].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6812_ (.D(_0995_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[14].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6813_ (.D(_0996_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[15].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6814_ (.D(_0997_),
    .GATE_N(net295),
    .Q(\stage_gen[3].mux_gen[15].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6815_ (.D(_0998_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[15].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6816_ (.D(_0999_),
    .GATE_N(net389),
    .Q(\stage_gen[3].mux_gen[15].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6817_ (.D(_1000_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[15].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6818_ (.D(_1001_),
    .GATE_N(net388),
    .Q(\stage_gen[3].mux_gen[16].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6819_ (.D(_1002_),
    .GATE_N(net296),
    .Q(\stage_gen[3].mux_gen[16].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6820_ (.D(_1003_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[16].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6821_ (.D(_1004_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[16].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6822_ (.D(_1005_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[16].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6823_ (.D(_1006_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[17].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6824_ (.D(_1007_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[17].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6825_ (.D(_1008_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[17].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6826_ (.D(_1009_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[17].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6827_ (.D(_1010_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[17].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6828_ (.D(_1011_),
    .GATE_N(net390),
    .Q(\stage_gen[3].mux_gen[18].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6829_ (.D(_1012_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[18].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6830_ (.D(_1013_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[18].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6831_ (.D(_1014_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[18].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6832_ (.D(_1015_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[18].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6833_ (.D(_1016_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[19].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6834_ (.D(_1017_),
    .GATE_N(net298),
    .Q(\stage_gen[3].mux_gen[19].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6835_ (.D(_1018_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[19].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6836_ (.D(_1019_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[19].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6837_ (.D(_1020_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[19].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6838_ (.D(_1026_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[20].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6839_ (.D(_1027_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[20].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6840_ (.D(_1028_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[20].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6841_ (.D(_1029_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[20].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6842_ (.D(_1030_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[20].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6843_ (.D(_1031_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[21].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6844_ (.D(_1032_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[21].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6845_ (.D(_1033_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[21].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6846_ (.D(_1034_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[21].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6847_ (.D(_1035_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[21].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6848_ (.D(_1036_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[22].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6849_ (.D(_1037_),
    .GATE_N(net297),
    .Q(\stage_gen[3].mux_gen[22].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6850_ (.D(_1038_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[22].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6851_ (.D(_1039_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[22].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6852_ (.D(_1040_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[22].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6853_ (.D(_1041_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[23].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6854_ (.D(_1042_),
    .GATE_N(net298),
    .Q(\stage_gen[3].mux_gen[23].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6855_ (.D(_1043_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[23].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6856_ (.D(_1044_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[23].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6857_ (.D(_1045_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[23].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6858_ (.D(_1046_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[24].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6859_ (.D(_1047_),
    .GATE_N(net298),
    .Q(\stage_gen[3].mux_gen[24].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6860_ (.D(_1048_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[24].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6861_ (.D(_1049_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[24].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6862_ (.D(_1050_),
    .GATE_N(net303),
    .Q(\stage_gen[3].mux_gen[24].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6863_ (.D(_1051_),
    .GATE_N(net391),
    .Q(\stage_gen[3].mux_gen[25].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6864_ (.D(_1052_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[25].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6865_ (.D(_1053_),
    .GATE_N(net400),
    .Q(\stage_gen[3].mux_gen[25].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6866_ (.D(_1054_),
    .GATE_N(net401),
    .Q(\stage_gen[3].mux_gen[25].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6867_ (.D(_1055_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[25].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6868_ (.D(_1056_),
    .GATE_N(net392),
    .Q(\stage_gen[3].mux_gen[26].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6869_ (.D(_1057_),
    .GATE_N(net298),
    .Q(\stage_gen[3].mux_gen[26].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6870_ (.D(_1058_),
    .GATE_N(net399),
    .Q(\stage_gen[3].mux_gen[26].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6871_ (.D(_1059_),
    .GATE_N(net398),
    .Q(\stage_gen[3].mux_gen[26].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6872_ (.D(_1060_),
    .GATE_N(net302),
    .Q(\stage_gen[3].mux_gen[26].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6873_ (.D(_1061_),
    .GATE_N(net397),
    .Q(\stage_gen[3].mux_gen[27].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6874_ (.D(_1062_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[27].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6875_ (.D(_1063_),
    .GATE_N(net401),
    .Q(\stage_gen[3].mux_gen[27].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6876_ (.D(_1064_),
    .GATE_N(net401),
    .Q(\stage_gen[3].mux_gen[27].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6877_ (.D(_1065_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[27].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6878_ (.D(_1066_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[28].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6879_ (.D(_1067_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[28].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6880_ (.D(_1068_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[28].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6881_ (.D(_1069_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[28].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6882_ (.D(_1070_),
    .GATE_N(net301),
    .Q(\stage_gen[3].mux_gen[28].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6883_ (.D(_1071_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[29].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6884_ (.D(_1072_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[29].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6885_ (.D(_1073_),
    .GATE_N(net397),
    .Q(\stage_gen[3].mux_gen[29].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6886_ (.D(_1074_),
    .GATE_N(net397),
    .Q(\stage_gen[3].mux_gen[29].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6887_ (.D(_1075_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[29].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6888_ (.D(_1081_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[30].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6889_ (.D(_1082_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[30].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6890_ (.D(_1083_),
    .GATE_N(net397),
    .Q(\stage_gen[3].mux_gen[30].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6891_ (.D(_1084_),
    .GATE_N(net394),
    .Q(\stage_gen[3].mux_gen[30].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6892_ (.D(_1085_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[30].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6893_ (.D(_1086_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[31].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6894_ (.D(_1087_),
    .GATE_N(net300),
    .Q(\stage_gen[3].mux_gen[31].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6895_ (.D(_1088_),
    .GATE_N(net397),
    .Q(\stage_gen[3].mux_gen[31].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6896_ (.D(_1089_),
    .GATE_N(net396),
    .Q(\stage_gen[3].mux_gen[31].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6897_ (.D(_1090_),
    .GATE_N(net299),
    .Q(\stage_gen[3].mux_gen[31].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_1324_),
    .Q(\stage_gen[4].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(clknet_3_5__leaf_CLK),
    .D(net514),
    .Q(\stage_gen[4].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(clknet_3_5__leaf_CLK),
    .D(net515),
    .Q(\stage_gen[4].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(clknet_3_5__leaf_CLK),
    .D(net506),
    .Q(\stage_gen[4].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net494),
    .Q(\stage_gen[4].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(clknet_3_5__leaf_CLK),
    .D(net507),
    .Q(\stage_gen[4].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(clknet_3_4__leaf_CLK),
    .D(net481),
    .Q(\stage_gen[4].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net508),
    .Q(\stage_gen[4].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(clknet_3_1__leaf_CLK),
    .D(net482),
    .Q(\stage_gen[4].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(clknet_3_4__leaf_CLK),
    .D(net484),
    .Q(\stage_gen[4].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_1334_),
    .Q(\stage_gen[4].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _6909_ (.D(_1126_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6910_ (.D(_1127_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6911_ (.D(_1128_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6912_ (.D(_1129_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6913_ (.D(_1130_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6914_ (.D(_1163_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6915_ (.D(_1164_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6916_ (.D(_1165_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6917_ (.D(_1166_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6918_ (.D(_1167_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6919_ (.D(_1168_),
    .GATE_N(net382),
    .Q(\stage_gen[4].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6920_ (.D(_1169_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6921_ (.D(_1170_),
    .GATE_N(net382),
    .Q(\stage_gen[4].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6922_ (.D(_1171_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6923_ (.D(_1172_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6924_ (.D(_1173_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6925_ (.D(_1174_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6926_ (.D(_1175_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6927_ (.D(_1176_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6928_ (.D(_1177_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6929_ (.D(_1178_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[4].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6930_ (.D(_1179_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[4].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6931_ (.D(_1180_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[4].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6932_ (.D(_1181_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[4].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6933_ (.D(_1182_),
    .GATE_N(net380),
    .Q(\stage_gen[4].mux_gen[4].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6934_ (.D(_1183_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[5].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6935_ (.D(_1184_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[5].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6936_ (.D(_1185_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[5].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6937_ (.D(_1186_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[5].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6938_ (.D(_1187_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[5].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6939_ (.D(_1188_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[6].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6940_ (.D(_1189_),
    .GATE_N(net380),
    .Q(\stage_gen[4].mux_gen[6].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6941_ (.D(_1190_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[6].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6942_ (.D(_1191_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[6].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6943_ (.D(_1192_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[6].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6944_ (.D(_1193_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[7].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6945_ (.D(_1194_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[7].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6946_ (.D(_1195_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[7].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6947_ (.D(_1196_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[7].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6948_ (.D(_1197_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[7].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6949_ (.D(_1198_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[8].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6950_ (.D(_1199_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[8].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6951_ (.D(_1200_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[8].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6952_ (.D(_1201_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[8].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6953_ (.D(_1202_),
    .GATE_N(net380),
    .Q(\stage_gen[4].mux_gen[8].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6954_ (.D(_1203_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[9].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6955_ (.D(_1204_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[9].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6956_ (.D(_1205_),
    .GATE_N(net387),
    .Q(\stage_gen[4].mux_gen[9].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6957_ (.D(_1206_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[9].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6958_ (.D(_1207_),
    .GATE_N(net378),
    .Q(\stage_gen[4].mux_gen[9].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6959_ (.D(_1133_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[10].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6960_ (.D(_1134_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[10].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6961_ (.D(_1135_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[10].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6962_ (.D(_1136_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[10].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6963_ (.D(_1137_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[10].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6964_ (.D(_1138_),
    .GATE_N(net384),
    .Q(\stage_gen[4].mux_gen[11].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6965_ (.D(_1139_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[11].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6966_ (.D(_1140_),
    .GATE_N(net387),
    .Q(\stage_gen[4].mux_gen[11].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6967_ (.D(_1141_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[11].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6968_ (.D(_1142_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[11].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6969_ (.D(_1143_),
    .GATE_N(net385),
    .Q(\stage_gen[4].mux_gen[12].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6970_ (.D(_1144_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[12].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6971_ (.D(_1145_),
    .GATE_N(net386),
    .Q(\stage_gen[4].mux_gen[12].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6972_ (.D(_1146_),
    .GATE_N(net387),
    .Q(\stage_gen[4].mux_gen[12].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6973_ (.D(_1147_),
    .GATE_N(net379),
    .Q(\stage_gen[4].mux_gen[12].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6974_ (.D(_1148_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[13].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6975_ (.D(_1149_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[13].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6976_ (.D(_1150_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[13].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6977_ (.D(_1151_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[13].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6978_ (.D(_1152_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[13].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6979_ (.D(_1153_),
    .GATE_N(net383),
    .Q(\stage_gen[4].mux_gen[14].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6980_ (.D(_1154_),
    .GATE_N(net377),
    .Q(\stage_gen[4].mux_gen[14].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6981_ (.D(_1155_),
    .GATE_N(net382),
    .Q(\stage_gen[4].mux_gen[14].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6982_ (.D(_1156_),
    .GATE_N(net382),
    .Q(\stage_gen[4].mux_gen[14].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6983_ (.D(_1157_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[14].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _6984_ (.D(_1158_),
    .GATE_N(net382),
    .Q(\stage_gen[4].mux_gen[15].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _6985_ (.D(_1159_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[15].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _6986_ (.D(_1160_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[15].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _6987_ (.D(_1161_),
    .GATE_N(net381),
    .Q(\stage_gen[4].mux_gen[15].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _6988_ (.D(_1162_),
    .GATE_N(net376),
    .Q(\stage_gen[4].mux_gen[15].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_1335_),
    .Q(\stage_gen[5].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_1336_),
    .Q(\stage_gen[5].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net485),
    .Q(\stage_gen[5].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net486),
    .Q(\stage_gen[5].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net487),
    .Q(\stage_gen[5].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net474),
    .Q(\stage_gen[5].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net463),
    .Q(\stage_gen[5].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net475),
    .Q(\stage_gen[5].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(clknet_3_7__leaf_CLK),
    .D(net464),
    .Q(\stage_gen[5].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net465),
    .Q(\stage_gen[5].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6999_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_1345_),
    .Q(\stage_gen[5].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _7000_ (.D(_1208_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7001_ (.D(_1209_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7002_ (.D(_1210_),
    .GATE_N(net440),
    .Q(\stage_gen[5].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7003_ (.D(_1211_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7004_ (.D(_1212_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7005_ (.D(_1215_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7006_ (.D(_1216_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7007_ (.D(_1217_),
    .GATE_N(net440),
    .Q(\stage_gen[5].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7008_ (.D(_1218_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7009_ (.D(_1219_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7010_ (.D(_1220_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7011_ (.D(_1221_),
    .GATE_N(net436),
    .Q(\stage_gen[5].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7012_ (.D(_1222_),
    .GATE_N(net440),
    .Q(\stage_gen[5].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7013_ (.D(_1223_),
    .GATE_N(net439),
    .Q(\stage_gen[5].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7014_ (.D(_1224_),
    .GATE_N(net436),
    .Q(\stage_gen[5].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7015_ (.D(_1225_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7016_ (.D(_1226_),
    .GATE_N(net436),
    .Q(\stage_gen[5].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7017_ (.D(_1227_),
    .GATE_N(net439),
    .Q(\stage_gen[5].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7018_ (.D(_1228_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7019_ (.D(_1229_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7020_ (.D(_1230_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[4].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7021_ (.D(_1231_),
    .GATE_N(net436),
    .Q(\stage_gen[5].mux_gen[4].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7022_ (.D(_1232_),
    .GATE_N(net439),
    .Q(\stage_gen[5].mux_gen[4].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7023_ (.D(_1233_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[4].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7024_ (.D(_1234_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[4].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7025_ (.D(_1235_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[5].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7026_ (.D(_1236_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[5].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7027_ (.D(_1237_),
    .GATE_N(net439),
    .Q(\stage_gen[5].mux_gen[5].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7028_ (.D(_1238_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[5].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7029_ (.D(_1239_),
    .GATE_N(net434),
    .Q(\stage_gen[5].mux_gen[5].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7030_ (.D(_1240_),
    .GATE_N(net438),
    .Q(\stage_gen[5].mux_gen[6].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7031_ (.D(_1241_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[6].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7032_ (.D(_1242_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[6].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7033_ (.D(_1243_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[6].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7034_ (.D(_1244_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[6].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7035_ (.D(_1245_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[7].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7036_ (.D(_1246_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[7].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7037_ (.D(_1247_),
    .GATE_N(net440),
    .Q(\stage_gen[5].mux_gen[7].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7038_ (.D(_1248_),
    .GATE_N(net437),
    .Q(\stage_gen[5].mux_gen[7].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7039_ (.D(_1249_),
    .GATE_N(net435),
    .Q(\stage_gen[5].mux_gen[7].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_1346_),
    .Q(\stage_gen[6].genblk1.clks.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7041_ (.CLK(clknet_3_2__leaf_CLK),
    .D(net495),
    .Q(\stage_gen[6].genblk1.clks.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net496),
    .Q(\stage_gen[6].genblk1.clks.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net476),
    .Q(\stage_gen[6].genblk1.clks.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7044_ (.CLK(clknet_3_6__leaf_CLK),
    .D(net466),
    .Q(\stage_gen[6].genblk1.clks.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7045_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net477),
    .Q(\stage_gen[6].genblk1.clks.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net467),
    .Q(\stage_gen[6].genblk1.clks.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7047_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net478),
    .Q(\stage_gen[6].genblk1.clks.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7048_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net497),
    .Q(\stage_gen[6].genblk1.clks.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7049_ (.CLK(clknet_3_3__leaf_CLK),
    .D(net498),
    .Q(\stage_gen[6].genblk1.clks.counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_1356_),
    .Q(\stage_gen[6].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _7051_ (.D(_1250_),
    .GATE_N(net433),
    .Q(\stage_gen[6].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7052_ (.D(_1251_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7053_ (.D(_1252_),
    .GATE_N(net433),
    .Q(\stage_gen[6].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7054_ (.D(_1253_),
    .GATE_N(_1255_),
    .Q(\stage_gen[6].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7055_ (.D(_1254_),
    .GATE_N(_1256_),
    .Q(\stage_gen[6].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7056_ (.D(_1257_),
    .GATE_N(net433),
    .Q(\stage_gen[6].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7057_ (.D(_1258_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7058_ (.D(_1259_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7059_ (.D(_1260_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7060_ (.D(_1261_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7061_ (.D(_1262_),
    .GATE_N(net433),
    .Q(\stage_gen[6].mux_gen[2].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7062_ (.D(_1263_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[2].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7063_ (.D(_1264_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[2].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7064_ (.D(_1265_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[2].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7065_ (.D(_1266_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[2].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7066_ (.D(_1267_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[3].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7067_ (.D(_1268_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[3].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7068_ (.D(_1269_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[3].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7069_ (.D(_1270_),
    .GATE_N(net432),
    .Q(\stage_gen[6].mux_gen[3].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7070_ (.D(_1271_),
    .GATE_N(net431),
    .Q(\stage_gen[6].mux_gen[3].S.IN1_L5 ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_1357_),
    .Q(\stage_gen[7].genblk1.clks.clk_o ));
 sky130_fd_sc_hd__dlxtn_1 _7072_ (.D(_1272_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7073_ (.D(_1273_),
    .GATE_N(_1278_),
    .Q(\stage_gen[7].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7074_ (.D(_1274_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7075_ (.D(_1275_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7076_ (.D(_1276_),
    .GATE_N(_1278_),
    .Q(\stage_gen[7].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7077_ (.D(_1279_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[1].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7078_ (.D(_1280_),
    .GATE_N(_1278_),
    .Q(\stage_gen[7].mux_gen[1].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7079_ (.D(_1281_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[1].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7080_ (.D(_1282_),
    .GATE_N(_1277_),
    .Q(\stage_gen[7].mux_gen[1].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7081_ (.D(_1283_),
    .GATE_N(_1278_),
    .Q(\stage_gen[7].mux_gen[1].S.IN1_L5 ));
 sky130_fd_sc_hd__dlxtn_1 _7082_ (.D(_1284_),
    .GATE_N(net455),
    .Q(\stage_gen[8].mux_gen[0].S.IN1_L1 ));
 sky130_fd_sc_hd__dlxtn_1 _7083_ (.D(_1285_),
    .GATE_N(clknet_1_1__leaf__1290_),
    .Q(\stage_gen[8].mux_gen[0].S.IN1_L2 ));
 sky130_fd_sc_hd__dlxtn_1 _7084_ (.D(clknet_1_0__leaf__1286_),
    .GATE_N(net454),
    .Q(\stage_gen[8].mux_gen[0].S.IN1_L3 ));
 sky130_fd_sc_hd__dlxtn_1 _7085_ (.D(_1287_),
    .GATE_N(net453),
    .Q(\stage_gen[8].mux_gen[0].S.IN1_L4 ));
 sky130_fd_sc_hd__dlxtn_1 _7086_ (.D(_1288_),
    .GATE_N(clknet_1_1__leaf__1290_),
    .Q(\stage_gen[8].mux_gen[0].S.IN1_L5 ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1286_ (.A(_1286_),
    .X(clknet_0__1286_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1290_ (.A(_1290_),
    .X(clknet_0__1290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2017_ (.A(_2017_),
    .X(clknet_0__2017_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2018_ (.A(_2018_),
    .X(clknet_0__2018_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2022_ (.A(_2022_),
    .X(clknet_0__2022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2023_ (.A(_2023_),
    .X(clknet_0__2023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2236_ (.A(_2236_),
    .X(clknet_0__2236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2678_ (.A(_2678_),
    .X(clknet_0__2678_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2681_ (.A(_2681_),
    .X(clknet_0__2681_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2683_ (.A(_2683_),
    .X(clknet_0__2683_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2684_ (.A(_2684_),
    .X(clknet_0__2684_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2695_ (.A(_2695_),
    .X(clknet_0__2695_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2703_ (.A(_2703_),
    .X(clknet_0__2703_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2706_ (.A(_2706_),
    .X(clknet_0__2706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2721_ (.A(_2721_),
    .X(clknet_0__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2724_ (.A(_2724_),
    .X(clknet_0__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2727_ (.A(_2727_),
    .X(clknet_0__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2730_ (.A(_2730_),
    .X(clknet_0__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2763_ (.A(_2763_),
    .X(clknet_0__2763_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2766_ (.A(_2766_),
    .X(clknet_0__2766_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2768_ (.A(_2768_),
    .X(clknet_0__2768_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2800_ (.A(_2800_),
    .X(clknet_0__2800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2803_ (.A(_2803_),
    .X(clknet_0__2803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2805_ (.A(_2805_),
    .X(clknet_0__2805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2830_ (.A(_2830_),
    .X(clknet_0__2830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2858_ (.A(_2858_),
    .X(clknet_0__2858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1286_ (.A(clknet_0__1286_),
    .X(clknet_1_0__leaf__1286_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1290_ (.A(clknet_0__1290_),
    .X(clknet_1_0__leaf__1290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2017_ (.A(clknet_0__2017_),
    .X(clknet_1_0__leaf__2017_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2018_ (.A(clknet_0__2018_),
    .X(clknet_1_0__leaf__2018_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2022_ (.A(clknet_0__2022_),
    .X(clknet_1_0__leaf__2022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2023_ (.A(clknet_0__2023_),
    .X(clknet_1_0__leaf__2023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2236_ (.A(clknet_0__2236_),
    .X(clknet_1_0__leaf__2236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2678_ (.A(clknet_0__2678_),
    .X(clknet_1_0__leaf__2678_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2681_ (.A(clknet_0__2681_),
    .X(clknet_1_0__leaf__2681_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2683_ (.A(clknet_0__2683_),
    .X(clknet_1_0__leaf__2683_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2684_ (.A(clknet_0__2684_),
    .X(clknet_1_0__leaf__2684_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2695_ (.A(clknet_0__2695_),
    .X(clknet_1_0__leaf__2695_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2703_ (.A(clknet_0__2703_),
    .X(clknet_1_0__leaf__2703_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2706_ (.A(clknet_0__2706_),
    .X(clknet_1_0__leaf__2706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2721_ (.A(clknet_0__2721_),
    .X(clknet_1_0__leaf__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2724_ (.A(clknet_0__2724_),
    .X(clknet_1_0__leaf__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2727_ (.A(clknet_0__2727_),
    .X(clknet_1_0__leaf__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2730_ (.A(clknet_0__2730_),
    .X(clknet_1_0__leaf__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2763_ (.A(clknet_0__2763_),
    .X(clknet_1_0__leaf__2763_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2766_ (.A(clknet_0__2766_),
    .X(clknet_1_0__leaf__2766_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2768_ (.A(clknet_0__2768_),
    .X(clknet_1_0__leaf__2768_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2800_ (.A(clknet_0__2800_),
    .X(clknet_1_0__leaf__2800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2803_ (.A(clknet_0__2803_),
    .X(clknet_1_0__leaf__2803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2805_ (.A(clknet_0__2805_),
    .X(clknet_1_0__leaf__2805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2830_ (.A(clknet_0__2830_),
    .X(clknet_1_0__leaf__2830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2858_ (.A(clknet_0__2858_),
    .X(clknet_1_0__leaf__2858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1286_ (.A(clknet_0__1286_),
    .X(clknet_1_1__leaf__1286_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1290_ (.A(clknet_0__1290_),
    .X(clknet_1_1__leaf__1290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2017_ (.A(clknet_0__2017_),
    .X(clknet_1_1__leaf__2017_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2018_ (.A(clknet_0__2018_),
    .X(clknet_1_1__leaf__2018_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2022_ (.A(clknet_0__2022_),
    .X(clknet_1_1__leaf__2022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2023_ (.A(clknet_0__2023_),
    .X(clknet_1_1__leaf__2023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2236_ (.A(clknet_0__2236_),
    .X(clknet_1_1__leaf__2236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2678_ (.A(clknet_0__2678_),
    .X(clknet_1_1__leaf__2678_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2681_ (.A(clknet_0__2681_),
    .X(clknet_1_1__leaf__2681_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2683_ (.A(clknet_0__2683_),
    .X(clknet_1_1__leaf__2683_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2684_ (.A(clknet_0__2684_),
    .X(clknet_1_1__leaf__2684_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2695_ (.A(clknet_0__2695_),
    .X(clknet_1_1__leaf__2695_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2703_ (.A(clknet_0__2703_),
    .X(clknet_1_1__leaf__2703_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2706_ (.A(clknet_0__2706_),
    .X(clknet_1_1__leaf__2706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2721_ (.A(clknet_0__2721_),
    .X(clknet_1_1__leaf__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2724_ (.A(clknet_0__2724_),
    .X(clknet_1_1__leaf__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2727_ (.A(clknet_0__2727_),
    .X(clknet_1_1__leaf__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2730_ (.A(clknet_0__2730_),
    .X(clknet_1_1__leaf__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2763_ (.A(clknet_0__2763_),
    .X(clknet_1_1__leaf__2763_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2766_ (.A(clknet_0__2766_),
    .X(clknet_1_1__leaf__2766_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2768_ (.A(clknet_0__2768_),
    .X(clknet_1_1__leaf__2768_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2800_ (.A(clknet_0__2800_),
    .X(clknet_1_1__leaf__2800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2803_ (.A(clknet_0__2803_),
    .X(clknet_1_1__leaf__2803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2805_ (.A(clknet_0__2805_),
    .X(clknet_1_1__leaf__2805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2830_ (.A(clknet_0__2830_),
    .X(clknet_1_1__leaf__2830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2858_ (.A(clknet_0__2858_),
    .X(clknet_1_1__leaf__2858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_2__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_3__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_4__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_5__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_6__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_7__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_2 fanout260 (.A(net264),
    .X(net260));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(net263),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 fanout264 (.A(net294),
    .X(net264));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(net267),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 fanout267 (.A(net272),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(net272),
    .X(net268));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout269 (.A(net272),
    .X(net269));
 sky130_fd_sc_hd__buf_2 fanout270 (.A(net272),
    .X(net270));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout272 (.A(net294),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_2 fanout274 (.A(net278),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(net278),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_2 fanout278 (.A(net294),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(net283),
    .X(net279));
 sky130_fd_sc_hd__buf_2 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(net294),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net288),
    .X(net284));
 sky130_fd_sc_hd__buf_2 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 fanout286 (.A(net288),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_2 fanout288 (.A(net293),
    .X(net288));
 sky130_fd_sc_hd__buf_2 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_2 fanout290 (.A(net292),
    .X(net290));
 sky130_fd_sc_hd__buf_2 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_2 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(_0006_),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_2 fanout296 (.A(net303),
    .X(net296));
 sky130_fd_sc_hd__buf_2 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout298 (.A(net303),
    .X(net298));
 sky130_fd_sc_hd__buf_2 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_2 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(net303),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(_0970_),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net315),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(net315),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(net315),
    .X(net306));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout307 (.A(net315),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net314),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 fanout309 (.A(net314),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net314),
    .X(net310));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout311 (.A(net314),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_2 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_2 fanout315 (.A(_0648_),
    .X(net315));
 sky130_fd_sc_hd__buf_2 fanout316 (.A(net321),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(net319),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__buf_2 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 fanout322 (.A(_0648_),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(net342),
    .X(net324));
 sky130_fd_sc_hd__buf_2 fanout325 (.A(net342),
    .X(net325));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout326 (.A(net342),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(net331),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(net331),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(net342),
    .X(net331));
 sky130_fd_sc_hd__buf_2 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_2 fanout333 (.A(net342),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 fanout334 (.A(net336),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 fanout336 (.A(net342),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 fanout337 (.A(net339),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_2 fanout339 (.A(net342),
    .X(net339));
 sky130_fd_sc_hd__buf_2 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 fanout342 (.A(_0005_),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net346),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 fanout344 (.A(net346),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_2 fanout347 (.A(net358),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net352),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(net358),
    .X(net352));
 sky130_fd_sc_hd__buf_2 fanout353 (.A(net355),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net358),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(_0005_),
    .X(net358));
 sky130_fd_sc_hd__buf_2 fanout359 (.A(net362),
    .X(net359));
 sky130_fd_sc_hd__buf_2 fanout360 (.A(net362),
    .X(net360));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 fanout362 (.A(net374),
    .X(net362));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(net374),
    .X(net365));
 sky130_fd_sc_hd__buf_2 fanout366 (.A(net370),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout370 (.A(net374),
    .X(net370));
 sky130_fd_sc_hd__buf_2 fanout371 (.A(net373),
    .X(net371));
 sky130_fd_sc_hd__buf_2 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(_0005_),
    .X(net375));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 fanout377 (.A(_1132_),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(net380),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 fanout380 (.A(_1132_),
    .X(net380));
 sky130_fd_sc_hd__buf_2 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 fanout383 (.A(net387),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 fanout384 (.A(net386),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(_1131_),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 fanout388 (.A(net393),
    .X(net388));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(net393),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_2 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout393 (.A(net402),
    .X(net393));
 sky130_fd_sc_hd__buf_2 fanout394 (.A(net402),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_2 fanout395 (.A(net402),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(net402),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(net401),
    .X(net399));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 fanout402 (.A(_0969_),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_4 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 fanout406 (.A(net409),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(_0647_),
    .X(net409));
 sky130_fd_sc_hd__buf_2 fanout410 (.A(net412),
    .X(net410));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net419),
    .X(net412));
 sky130_fd_sc_hd__buf_2 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout414 (.A(net419),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(net419),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(net418),
    .X(net416));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_2 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(_0647_),
    .X(net419));
 sky130_fd_sc_hd__buf_2 fanout420 (.A(net430),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(net430),
    .X(net421));
 sky130_fd_sc_hd__buf_2 fanout422 (.A(net428),
    .X(net422));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout423 (.A(net428),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(net428),
    .X(net424));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout425 (.A(net428),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(net428),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(net430),
    .X(net428));
 sky130_fd_sc_hd__buf_2 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(_0647_),
    .X(net430));
 sky130_fd_sc_hd__buf_2 fanout431 (.A(_1256_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(_1255_),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 fanout434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(_1214_),
    .X(net435));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout436 (.A(_1214_),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net440),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_2 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 fanout440 (.A(_1213_),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(PAR_IN[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(PAR_IN[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(PAR_IN[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(PAR_IN[190]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(PAR_IN[191]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(PAR_IN[192]),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 input104 (.A(PAR_IN[193]),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(PAR_IN[194]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(PAR_IN[195]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(PAR_IN[196]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(PAR_IN[197]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(PAR_IN[198]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(PAR_IN[109]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(PAR_IN[199]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(PAR_IN[19]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(PAR_IN[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(PAR_IN[200]),
    .X(net113));
 sky130_fd_sc_hd__dlymetal6s2s_1 input114 (.A(PAR_IN[201]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(PAR_IN[202]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(PAR_IN[203]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(PAR_IN[204]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(PAR_IN[205]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(PAR_IN[206]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(PAR_IN[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(PAR_IN[207]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(PAR_IN[208]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(PAR_IN[209]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(PAR_IN[20]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(PAR_IN[210]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(PAR_IN[211]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(PAR_IN[212]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(PAR_IN[213]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(PAR_IN[214]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(PAR_IN[215]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(PAR_IN[110]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(PAR_IN[216]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(PAR_IN[217]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(PAR_IN[218]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(PAR_IN[219]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(PAR_IN[21]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(PAR_IN[220]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(PAR_IN[221]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(PAR_IN[222]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(PAR_IN[223]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(PAR_IN[224]),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(PAR_IN[111]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(PAR_IN[225]),
    .X(net140));
 sky130_fd_sc_hd__buf_2 input141 (.A(PAR_IN[226]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(PAR_IN[227]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(PAR_IN[228]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(PAR_IN[229]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(PAR_IN[22]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(PAR_IN[230]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(PAR_IN[231]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(PAR_IN[232]),
    .X(net148));
 sky130_fd_sc_hd__dlymetal6s2s_1 input149 (.A(PAR_IN[233]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(PAR_IN[112]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(PAR_IN[234]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(PAR_IN[235]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(PAR_IN[236]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(PAR_IN[237]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(PAR_IN[238]),
    .X(net154));
 sky130_fd_sc_hd__buf_2 input155 (.A(PAR_IN[239]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(PAR_IN[23]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(PAR_IN[240]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(PAR_IN[241]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(PAR_IN[242]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(PAR_IN[113]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(PAR_IN[243]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(PAR_IN[244]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(PAR_IN[245]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(PAR_IN[246]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(PAR_IN[247]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(PAR_IN[248]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(PAR_IN[249]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 input167 (.A(PAR_IN[24]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(PAR_IN[250]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(PAR_IN[251]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(PAR_IN[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(PAR_IN[252]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(PAR_IN[253]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(PAR_IN[254]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(PAR_IN[255]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(PAR_IN[25]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(PAR_IN[26]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 input176 (.A(PAR_IN[27]),
    .X(net176));
 sky130_fd_sc_hd__buf_2 input177 (.A(PAR_IN[28]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(PAR_IN[29]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(PAR_IN[2]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(PAR_IN[115]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input180 (.A(PAR_IN[30]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(PAR_IN[31]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 input182 (.A(PAR_IN[32]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(PAR_IN[33]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(PAR_IN[34]),
    .X(net184));
 sky130_fd_sc_hd__buf_2 input185 (.A(PAR_IN[35]),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 input186 (.A(PAR_IN[36]),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 input187 (.A(PAR_IN[37]),
    .X(net187));
 sky130_fd_sc_hd__buf_2 input188 (.A(PAR_IN[38]),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(PAR_IN[39]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(PAR_IN[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input190 (.A(PAR_IN[3]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(PAR_IN[40]),
    .X(net191));
 sky130_fd_sc_hd__buf_2 input192 (.A(PAR_IN[41]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(PAR_IN[42]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(PAR_IN[43]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(PAR_IN[44]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(PAR_IN[45]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input197 (.A(PAR_IN[46]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(PAR_IN[47]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(PAR_IN[48]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(PAR_IN[100]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(PAR_IN[117]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(PAR_IN[49]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(PAR_IN[4]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 input202 (.A(PAR_IN[50]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(PAR_IN[51]),
    .X(net203));
 sky130_fd_sc_hd__buf_2 input204 (.A(PAR_IN[52]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(PAR_IN[53]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(PAR_IN[54]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 input207 (.A(PAR_IN[55]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(PAR_IN[56]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(PAR_IN[57]),
    .X(net209));
 sky130_fd_sc_hd__buf_2 input21 (.A(PAR_IN[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(PAR_IN[58]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(PAR_IN[59]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(PAR_IN[5]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(PAR_IN[60]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(PAR_IN[61]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(PAR_IN[62]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(PAR_IN[63]),
    .X(net216));
 sky130_fd_sc_hd__buf_2 input217 (.A(PAR_IN[64]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 input218 (.A(PAR_IN[65]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 input219 (.A(PAR_IN[66]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(PAR_IN[119]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(PAR_IN[67]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(PAR_IN[68]),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(PAR_IN[69]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(PAR_IN[6]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(PAR_IN[70]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_4 input225 (.A(PAR_IN[71]),
    .X(net225));
 sky130_fd_sc_hd__buf_2 input226 (.A(PAR_IN[72]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 input227 (.A(PAR_IN[73]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(PAR_IN[74]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(PAR_IN[75]),
    .X(net229));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(PAR_IN[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(PAR_IN[76]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(PAR_IN[77]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(PAR_IN[78]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(PAR_IN[79]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 input234 (.A(PAR_IN[7]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(PAR_IN[80]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(PAR_IN[81]),
    .X(net236));
 sky130_fd_sc_hd__dlymetal6s2s_1 input237 (.A(PAR_IN[82]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(PAR_IN[83]),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input239 (.A(PAR_IN[84]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(PAR_IN[120]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(PAR_IN[85]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 input241 (.A(PAR_IN[86]),
    .X(net241));
 sky130_fd_sc_hd__buf_2 input242 (.A(PAR_IN[87]),
    .X(net242));
 sky130_fd_sc_hd__buf_2 input243 (.A(PAR_IN[88]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(PAR_IN[89]),
    .X(net244));
 sky130_fd_sc_hd__dlymetal6s2s_1 input245 (.A(PAR_IN[8]),
    .X(net245));
 sky130_fd_sc_hd__dlymetal6s2s_1 input246 (.A(PAR_IN[90]),
    .X(net246));
 sky130_fd_sc_hd__dlymetal6s2s_1 input247 (.A(PAR_IN[91]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 input248 (.A(PAR_IN[92]),
    .X(net248));
 sky130_fd_sc_hd__buf_2 input249 (.A(PAR_IN[93]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(PAR_IN[121]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input250 (.A(PAR_IN[94]),
    .X(net250));
 sky130_fd_sc_hd__buf_2 input251 (.A(PAR_IN[95]),
    .X(net251));
 sky130_fd_sc_hd__buf_2 input252 (.A(PAR_IN[96]),
    .X(net252));
 sky130_fd_sc_hd__dlymetal6s2s_1 input253 (.A(PAR_IN[97]),
    .X(net253));
 sky130_fd_sc_hd__dlymetal6s2s_1 input254 (.A(PAR_IN[98]),
    .X(net254));
 sky130_fd_sc_hd__buf_2 input255 (.A(PAR_IN[99]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 input256 (.A(PAR_IN[9]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(RESET),
    .X(net257));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(PAR_IN[122]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(PAR_IN[123]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(PAR_IN[124]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(PAR_IN[125]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(PAR_IN[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(PAR_IN[126]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(PAR_IN[127]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(PAR_IN[128]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(PAR_IN[129]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(PAR_IN[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(PAR_IN[130]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(PAR_IN[131]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(PAR_IN[132]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(PAR_IN[133]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(PAR_IN[134]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(PAR_IN[102]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(PAR_IN[135]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(PAR_IN[136]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(PAR_IN[137]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(PAR_IN[138]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(PAR_IN[139]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(PAR_IN[13]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(PAR_IN[140]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(PAR_IN[141]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(PAR_IN[142]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(PAR_IN[143]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(PAR_IN[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input50 (.A(PAR_IN[144]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(PAR_IN[145]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(PAR_IN[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(PAR_IN[147]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(PAR_IN[148]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(PAR_IN[149]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(PAR_IN[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(PAR_IN[150]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(PAR_IN[151]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(PAR_IN[152]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(PAR_IN[104]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(PAR_IN[153]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(PAR_IN[154]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(PAR_IN[155]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(PAR_IN[156]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(PAR_IN[157]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(PAR_IN[158]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(PAR_IN[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(PAR_IN[15]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(PAR_IN[160]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(PAR_IN[161]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(PAR_IN[105]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(PAR_IN[162]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(PAR_IN[163]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(PAR_IN[164]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(PAR_IN[165]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(PAR_IN[166]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(PAR_IN[167]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(PAR_IN[168]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(PAR_IN[169]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(PAR_IN[16]),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 input79 (.A(PAR_IN[170]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(PAR_IN[106]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(PAR_IN[171]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(PAR_IN[172]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(PAR_IN[173]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(PAR_IN[174]),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(PAR_IN[175]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(PAR_IN[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(PAR_IN[177]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(PAR_IN[178]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(PAR_IN[179]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(PAR_IN[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(PAR_IN[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(PAR_IN[180]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(PAR_IN[181]),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 input92 (.A(PAR_IN[182]),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input93 (.A(PAR_IN[183]),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(PAR_IN[184]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(PAR_IN[185]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(PAR_IN[186]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(PAR_IN[187]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(PAR_IN[188]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(PAR_IN[189]),
    .X(net99));
 sky130_fd_sc_hd__inv_2 net399_2 (.A(clknet_3_5__leaf_CLK),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 net399_3 (.A(clknet_3_7__leaf_CLK),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 net399_4 (.A(clknet_3_7__leaf_CLK),
    .Y(net444));
 sky130_fd_sc_hd__clkbuf_1 output258 (.A(net258),
    .X(SERIAL_OUT));
endmodule

